0,0
1,0
2,0
3,0
4,0
5,0
6,0
7,0
8,0
9,0
10,0
11,0
12,0
13,0
14,0
15,0
16,0
17,0
18,0
19,0
20,0
21,0
22,0
23,0
24,0
25,0
26,0
27,0
28,0
29,0
30,0
31,0
32,0
33,0
34,0
35,0
36,0
37,0
38,0
39,0
40,0
41,0
42,0
43,0
44,0
45,0
46,1
47,1
48,1
49,1
50,1
51,1
52,1
53,1
54,1
55,1
56,1
57,1
58,1
59,1
60,1
61,1
62,1
63,1
64,1
65,1
66,1
67,1
68,1
69,1
70,1
71,1
72,1
73,1
74,1
75,1
76,1
77,1
78,1
79,1
80,1
81,1
82,1
83,1
84,1
85,1
86,1
87,1
88,1
89,1
90,1
91,1
92,2
93,2
94,2
95,2
96,2
97,2
98,2
99,2
100,2
101,2
102,2
103,2
104,2
105,2
106,2
107,2
108,2
109,2
110,2
111,2
112,2
113,2
114,2
115,2
116,2
117,2
118,2
119,2
120,2
121,2
122,2
123,2
124,2
125,2
126,2
127,2
128,2
129,2
130,2
131,2
132,2
133,2
134,2
135,2
136,2
137,2
138,3
139,3
140,3
141,3
142,3
143,3
144,3
145,3
146,3
147,3
148,3
149,3
150,3
151,3
152,3
153,3
154,3
155,3
156,3
157,3
158,3
159,3
160,3
161,3
162,3
163,3
164,3
165,3
166,3
167,3
168,3
169,3
170,3
171,3
172,3
173,3
174,3
175,3
176,3
177,3
178,3
179,3
180,3
181,3
182,3
183,3
184,4
185,4
186,4
187,4
188,4
189,4
190,4
191,4
192,4
193,4
194,4
195,4
196,4
197,4
198,4
199,4
200,4
201,4
202,4
203,4
204,4
205,4
206,4
207,4
208,4
209,4
210,4
211,4
212,4
213,4
214,4
215,4
216,4
217,4
218,4
219,4
220,4
221,4
222,4
223,4
224,4
225,4
226,4
227,4
228,4
229,4
230,5
231,5
232,5
233,5
234,5
235,5
236,5
237,5
238,5
239,5
240,5
241,5
242,5
243,5
244,5
245,5
246,5
247,5
248,5
249,5
250,5
251,5
252,5
253,5
254,5
255,5
256,5
257,5
258,5
259,5
260,5
261,5
262,5
263,5
264,5
265,5
266,5
267,5
268,5
269,5
270,5
271,5
272,5
273,5
274,5
275,5
276,6
277,6
278,6
279,6
280,6
281,6
282,6
283,6
284,6
285,6
286,6
287,6
288,6
289,6
290,6
291,6
292,6
293,6
294,6
295,6
296,6
297,6
298,6
299,6
300,6
301,6
302,6
303,6
304,6
305,6
306,6
307,6
308,6
309,6
310,6
311,6
312,6
313,6
314,6
315,6
316,6
317,6
318,6
319,6
320,6
321,6
322,7
323,7
324,7
325,7
326,7
327,7
328,7
329,7
330,7
331,7
332,7
333,7
334,7
335,7
336,7
337,7
338,7
339,7
340,7
341,7
342,7
343,7
344,7
345,7
346,7
347,7
348,7
349,7
350,7
351,7
352,7
353,7
354,7
355,7
356,7
357,7
358,7
359,7
360,7
361,7
362,7
363,7
364,7
365,7
366,7
367,7
368,8
369,8
370,8
371,8
372,8
373,8
374,8
375,8
376,8
377,8
378,8
379,8
380,8
381,8
382,8
383,8
384,8
385,8
386,8
387,8
388,8
389,8
390,8
391,8
392,8
393,8
394,8
395,8
396,8
397,8
398,8
399,8
400,8
401,8
402,8
403,8
404,8
405,8
406,8
407,8
408,8
409,8
410,8
411,8
412,8
413,8
414,9
415,9
416,9
417,9
418,9
419,9
420,9
421,9
422,9
423,9
424,9
425,9
426,9
427,9
428,9
429,9
430,9
431,9
432,9
433,9
434,9
435,9
436,9
437,9
438,9
439,9
440,9
441,9
442,9
443,9
444,9
445,9
446,9
447,9
448,9
449,9
450,9
451,9
452,9
453,9
454,9
455,9
456,9
457,9
458,9
459,9
460,10
461,10
462,10
463,10
464,10
465,10
466,10
467,10
468,10
469,10
470,10
471,10
472,10
473,10
474,10
475,10
476,10
477,10
478,10
479,10
480,10
481,10
482,10
483,10
484,10
485,10
486,10
487,10
488,10
489,10
490,10
491,10
492,10
493,10
494,10
495,10
496,10
497,10
498,10
499,10
500,10
501,10
502,10
503,10
504,10
505,10
506,11
507,11
508,11
509,11
510,11
511,11
512,11
513,11
514,11
515,11
516,11
517,11
518,11
519,11
520,11
521,11
522,11
523,11
524,11
525,11
526,11
527,11
528,11
529,11
530,11
531,11
532,11
533,11
534,11
535,11
536,11
537,11
538,11
539,11
540,11
541,11
542,11
543,11
544,11
545,11
546,11
547,11
548,11
549,11
550,11
551,11
552,12
553,12
554,12
555,12
556,12
557,12
558,12
559,12
560,12
561,12
562,12
563,12
564,12
565,12
566,12
567,12
568,12
569,12
570,12
571,12
572,12
573,12
574,12
575,12
576,12
577,12
578,12
579,12
580,12
581,12
582,12
583,12
584,12
585,12
586,12
587,12
588,12
589,12
590,12
591,12
592,12
593,12
594,12
595,12
596,12
597,12
598,13
599,13
600,13
601,13
602,13
603,13
604,13
605,13
606,13
607,13
608,13
609,13
610,13
611,13
612,13
613,13
614,13
615,13
616,13
617,13
618,13
619,13
620,13
621,13
622,13
623,13
624,13
625,13
626,13
627,13
628,13
629,13
630,13
631,13
632,13
633,13
634,13
635,13
636,13
637,13
638,13
639,13
640,13
641,13
642,13
643,13
644,14
645,14
646,14
647,14
648,14
649,14
650,14
651,14
652,14
653,14
654,14
655,14
656,14
657,14
658,14
659,14
660,14
661,14
662,14
663,14
664,14
665,14
666,14
667,14
668,14
669,14
670,14
671,14
672,14
673,14
674,14
675,14
676,14
677,14
678,14
679,14
680,14
681,14
682,14
683,14
684,14
685,14
686,14
687,14
688,14
689,14
690,15
691,15
692,15
693,15
694,15
695,15
696,15
697,15
698,15
699,15
700,15
701,15
702,15
703,15
704,15
705,15
706,15
707,15
708,15
709,15
710,15
711,15
712,15
713,15
714,15
715,15
716,15
717,15
718,15
719,15
720,15
721,15
722,15
723,15
724,15
725,15
726,15
727,15
728,15
729,15
730,15
731,15
732,15
733,15
734,15
735,15
736,16
737,16
738,16
739,16
740,16
741,16
742,16
743,16
744,16
745,16
746,16
747,16
748,16
749,16
750,16
751,16
752,16
753,16
754,16
755,16
756,16
757,16
758,16
759,16
760,16
761,16
762,16
763,16
764,16
765,16
766,16
767,16
768,16
769,16
770,16
771,16
772,16
773,16
774,16
775,16
776,16
777,16
778,16
779,16
780,16
781,16
782,17
783,17
784,17
785,17
786,17
787,17
788,17
789,17
790,17
791,17
792,17
793,17
794,17
795,17
796,17
797,17
798,17
799,17
800,17
801,17
802,17
803,17
804,17
805,17
806,17
807,17
808,17
809,17
810,17
811,17
812,17
813,17
814,17
815,17
816,17
817,17
818,17
819,17
820,17
821,17
822,17
823,17
824,17
825,17
826,17
827,17
828,18
829,18
830,18
831,18
832,18
833,18
834,18
835,18
836,18
837,18
838,18
839,18
840,18
841,18
842,18
843,18
844,18
845,18
846,18
847,18
848,18
849,18
850,18
851,18
852,18
853,18
854,18
855,18
856,18
857,18
858,18
859,18
860,18
861,18
862,18
863,18
864,18
865,18
866,18
867,18
868,18
869,18
870,18
871,18
872,18
873,18
874,19
875,19
876,19
877,19
878,19
879,19
880,19
881,19
882,19
883,19
884,19
885,19
886,19
887,19
888,19
889,19
890,19
891,19
892,19
893,19
894,19
895,19
896,19
897,19
898,19
899,19
900,19
901,19
902,19
903,19
904,19
905,19
906,19
907,19
908,19
909,19
910,19
911,19
912,19
913,19
914,19
915,19
916,19
917,19
918,19
919,19
920,20
921,20
922,20
923,20
924,20
925,20
926,20
927,20
928,20
929,20
930,20
931,20
932,20
933,20
934,20
935,20
936,20
937,20
938,20
939,20
940,20
941,20
942,20
943,20
944,20
945,20
946,20
947,20
948,20
949,20
950,20
951,20
952,20
953,20
954,20
955,20
956,20
957,20
958,20
959,20
960,20
961,20
962,20
963,20
964,20
965,20
966,21
967,21
968,21
969,21
970,21
971,21
972,21
973,21
974,21
975,21
976,21
977,21
978,21
979,21
980,21
981,21
982,21
983,21
984,21
985,21
986,21
987,21
988,21
989,21
990,21
991,21
992,21
993,21
994,21
995,21
996,21
997,21
998,21
999,21
1000,21
1001,21
1002,21
1003,21
1004,21
1005,21
1006,21
1007,21
1008,21
1009,21
1010,21
1011,21
1012,22
1013,22
1014,22
1015,22
1016,22
1017,22
1018,22
1019,22
1020,22
1021,22
1022,22
1023,22
1024,22
1025,22
1026,22
1027,22
1028,22
1029,22
1030,22
1031,22
1032,22
1033,22
1034,22
1035,22
1036,22
1037,22
1038,22
1039,22
1040,22
1041,22
1042,22
1043,22
1044,22
1045,22
1046,22
1047,22
1048,22
1049,22
1050,22
1051,22
1052,22
1053,22
1054,22
1055,22
1056,22
1057,22
1058,23
1059,23
1060,23
1061,23
1062,23
1063,23
1064,23
1065,23
1066,23
1067,23
1068,23
1069,23
1070,23
1071,23
1072,23
1073,23
1074,23
1075,23
1076,23
1077,23
1078,23
1079,23
1080,23
1081,23
1082,23
1083,23
1084,23
1085,23
1086,23
1087,23
1088,23
1089,23
1090,23
1091,23
1092,23
1093,23
1094,23
1095,23
1096,23
1097,23
1098,23
1099,23
1100,23
1101,23
1102,23
1103,23
1104,24
1105,24
1106,24
1107,24
1108,24
1109,24
1110,24
1111,24
1112,24
1113,24
1114,24
1115,24
1116,24
1117,24
1118,24
1119,24
1120,24
1121,24
1122,24
1123,24
1124,24
1125,24
1126,24
1127,24
1128,24
1129,24
1130,24
1131,24
1132,24
1133,24
1134,24
1135,24
1136,24
1137,24
1138,24
1139,24
1140,24
1141,24
1142,24
1143,24
1144,24
1145,24
1146,24
1147,24
1148,24
1149,24
1150,25
1151,25
1152,25
1153,25
1154,25
1155,25
1156,25
1157,25
1158,25
1159,25
1160,25
1161,25
1162,25
1163,25
1164,25
1165,25
1166,25
1167,25
1168,25
1169,25
1170,25
1171,25
1172,25
1173,25
1174,25
1175,25
1176,25
1177,25
1178,25
1179,25
1180,25
1181,25
1182,25
1183,25
1184,25
1185,25
1186,25
1187,25
1188,25
1189,25
1190,25
1191,25
1192,25
1193,25
1194,25
1195,25
1196,26
1197,26
1198,26
1199,26
1200,26
1201,26
1202,26
1203,26
1204,26
1205,26
1206,26
1207,26
1208,26
1209,26
1210,26
1211,26
1212,26
1213,26
1214,26
1215,26
1216,26
1217,26
1218,26
1219,26
1220,26
1221,26
1222,26
1223,26
1224,26
1225,26
1226,26
1227,26
1228,26
1229,26
1230,26
1231,26
1232,26
1233,26
1234,26
1235,26
1236,26
1237,26
1238,26
1239,26
1240,26
1241,26
1242,27
1243,27
1244,27
1245,27
1246,27
1247,27
1248,27
1249,27
1250,27
1251,27
1252,27
1253,27
1254,27
1255,27
1256,27
1257,27
1258,27
1259,27
1260,27
1261,27
1262,27
1263,27
1264,27
1265,27
1266,27
1267,27
1268,27
1269,27
1270,27
1271,27
1272,27
1273,27
1274,27
1275,27
1276,27
1277,27
1278,27
1279,27
1280,27
1281,27
1282,27
1283,27
1284,27
1285,27
1286,27
1287,27
1288,28
1289,28
1290,28
1291,28
1292,28
1293,28
1294,28
1295,28
1296,28
1297,28
1298,28
1299,28
1300,28
1301,28
1302,28
1303,28
1304,28
1305,28
1306,28
1307,28
1308,28
1309,28
1310,28
1311,28
1312,28
1313,28
1314,28
1315,28
1316,28
1317,28
1318,28
1319,28
1320,28
1321,28
1322,28
1323,28
1324,28
1325,28
1326,28
1327,28
1328,28
1329,28
1330,28
1331,28
1332,28
1333,28
1334,29
1335,29
1336,29
1337,29
1338,29
1339,29
1340,29
1341,29
1342,29
1343,29
1344,29
1345,29
1346,29
1347,29
1348,29
1349,29
1350,29
1351,29
1352,29
1353,29
1354,29
1355,29
1356,29
1357,29
1358,29
1359,29
1360,29
1361,29
1362,29
1363,29
1364,29
1365,29
1366,29
1367,29
1368,29
1369,29
1370,29
1371,29
1372,29
1373,29
1374,29
1375,29
1376,29
1377,29
1378,29
1379,29
1380,30
1381,30
1382,30
1383,30
1384,30
1385,30
1386,30
1387,30
1388,30
1389,30
1390,30
1391,30
1392,30
1393,30
1394,30
1395,30
1396,30
1397,30
1398,30
1399,30
1400,30
1401,30
1402,30
1403,30
1404,30
1405,30
1406,30
1407,30
1408,30
1409,30
1410,30
1411,30
1412,30
1413,30
1414,30
1415,30
1416,30
1417,30
1418,30
1419,30
1420,30
1421,30
1422,30
1423,30
1424,30
1425,30
1426,31
1427,31
1428,31
1429,31
1430,31
1431,31
1432,31
1433,31
1434,31
1435,31
1436,31
1437,31
1438,31
1439,31
1440,31
1441,31
1442,31
1443,31
1444,31
1445,31
1446,31
1447,31
1448,31
1449,31
1450,31
1451,31
1452,31
1453,31
1454,31
1455,31
1456,31
1457,31
1458,31
1459,31
1460,31
1461,31
1462,31
1463,31
1464,31
1465,31
1466,31
1467,31
1468,31
1469,31
1470,31
1471,31
1472,32
1473,32
1474,32
1475,32
1476,32
1477,32
1478,32
1479,32
1480,32
1481,32
1482,32
1483,32
1484,32
1485,32
1486,32
1487,32
1488,32
1489,32
1490,32
1491,32
1492,32
1493,32
1494,32
1495,32
1496,32
1497,32
1498,32
1499,32
1500,32
1501,32
1502,32
1503,32
1504,32
1505,32
1506,32
1507,32
1508,32
1509,32
1510,32
1511,32
1512,32
1513,32
1514,32
1515,32
1516,32
1517,32
1518,33
1519,33
1520,33
1521,33
1522,33
1523,33
1524,33
1525,33
1526,33
1527,33
1528,33
1529,33
1530,33
1531,33
1532,33
1533,33
1534,33
1535,33
1536,33
1537,33
1538,33
1539,33
1540,33
1541,33
1542,33
1543,33
1544,33
1545,33
1546,33
1547,33
1548,33
1549,33
1550,33
1551,33
1552,33
1553,33
1554,33
1555,33
1556,33
1557,33
1558,33
1559,33
1560,33
1561,33
1562,33
1563,33
1564,34
1565,34
1566,34
1567,34
1568,34
1569,34
1570,34
1571,34
1572,34
1573,34
1574,34
1575,34
1576,34
1577,34
1578,34
1579,34
1580,34
1581,34
1582,34
1583,34
1584,34
1585,34
1586,34
1587,34
1588,34
1589,34
1590,34
1591,34
1592,34
1593,34
1594,34
1595,34
1596,34
1597,34
1598,34
1599,34
1600,34
1601,34
1602,34
1603,34
1604,34
1605,34
1606,34
1607,34
1608,34
1609,34
1610,35
1611,35
1612,35
1613,35
1614,35
1615,35
1616,35
1617,35
1618,35
1619,35
1620,35
1621,35
1622,35
1623,35
1624,35
1625,35
1626,35
1627,35
1628,35
1629,35
1630,35
1631,35
1632,35
1633,35
1634,35
1635,35
1636,35
1637,35
1638,35
1639,35
1640,35
1641,35
1642,35
1643,35
1644,35
1645,35
1646,35
1647,35
1648,35
1649,35
1650,35
1651,35
1652,35
1653,35
1654,35
1655,35
1656,36
1657,36
1658,36
1659,36
1660,36
1661,36
1662,36
1663,36
1664,36
1665,36
1666,36
1667,36
1668,36
1669,36
1670,36
1671,36
1672,36
1673,36
1674,36
1675,36
1676,36
1677,36
1678,36
1679,36
1680,36
1681,36
1682,36
1683,36
1684,36
1685,36
1686,36
1687,36
1688,36
1689,36
1690,36
1691,36
1692,36
1693,36
1694,36
1695,36
1696,36
1697,36
1698,36
1699,36
1700,36
1701,36
1702,37
1703,37
1704,37
1705,37
1706,37
1707,37
1708,37
1709,37
1710,37
1711,37
1712,37
1713,37
1714,37
1715,37
1716,37
1717,37
1718,37
1719,37
1720,37
1721,37
1722,37
1723,37
1724,37
1725,37
1726,37
1727,37
1728,37
1729,37
1730,37
1731,37
1732,37
1733,37
1734,37
1735,37
1736,37
1737,37
1738,37
1739,37
1740,37
1741,37
1742,37
1743,37
1744,37
1745,37
1746,37
1747,37
1748,38
1749,38
1750,38
1751,38
1752,38
1753,38
1754,38
1755,38
1756,38
1757,38
1758,38
1759,38
1760,38
1761,38
1762,38
1763,38
1764,38
1765,38
1766,38
1767,38
1768,38
1769,38
1770,38
1771,38
1772,38
1773,38
1774,38
1775,38
1776,38
1777,38
1778,38
1779,38
1780,38
1781,38
1782,38
1783,38
1784,38
1785,38
1786,38
1787,38
1788,38
1789,38
1790,38
1791,38
1792,38
1793,38
1794,39
1795,39
1796,39
1797,39
1798,39
1799,39
1800,39
1801,39
1802,39
1803,39
1804,39
1805,39
1806,39
1807,39
1808,39
1809,39
1810,39
1811,39
1812,39
1813,39
1814,39
1815,39
1816,39
1817,39
1818,39
1819,39
1820,39
1821,39
1822,39
1823,39
1824,39
1825,39
1826,39
1827,39
1828,39
1829,39
1830,39
1831,39
1832,39
1833,39
1834,39
1835,39
1836,39
1837,39
1838,39
1839,39
1840,40
1841,40
1842,40
1843,40
1844,40
1845,40
1846,40
1847,40
1848,40
1849,40
1850,40
1851,40
1852,40
1853,40
1854,40
1855,40
1856,40
1857,40
1858,40
1859,40
1860,40
1861,40
1862,40
1863,40
1864,40
1865,40
1866,40
1867,40
1868,40
1869,40
1870,40
1871,40
1872,40
1873,40
1874,40
1875,40
1876,40
1877,40
1878,40
1879,40
1880,40
1881,40
1882,40
1883,40
1884,40
1885,40
1886,41
1887,41
1888,41
1889,41
1890,41
1891,41
1892,41
1893,41
1894,41
1895,41
1896,41
1897,41
1898,41
1899,41
1900,41
1901,41
1902,41
1903,41
1904,41
1905,41
1906,41
1907,41
1908,41
1909,41
1910,41
1911,41
1912,41
1913,41
1914,41
1915,41
1916,41
1917,41
1918,41
1919,41
1920,41
1921,41
1922,41
1923,41
1924,41
1925,41
1926,41
1927,41
1928,41
1929,41
1930,41
1931,41
1932,42
1933,42
1934,42
1935,42
1936,42
1937,42
1938,42
1939,42
1940,42
1941,42
1942,42
1943,42
1944,42
1945,42
1946,42
1947,42
1948,42
1949,42
1950,42
1951,42
1952,42
1953,42
1954,42
1955,42
1956,42
1957,42
1958,42
1959,42
1960,42
1961,42
1962,42
1963,42
1964,42
1965,42
1966,42
1967,42
1968,42
1969,42
1970,42
1971,42
1972,42
1973,42
1974,42
1975,42
1976,42
1977,42
1978,43
1979,43
1980,43
1981,43
1982,43
1983,43
1984,43
1985,43
1986,43
1987,43
1988,43
1989,43
1990,43
1991,43
1992,43
1993,43
1994,43
1995,43
1996,43
1997,43
1998,43
1999,43
2000,43
2001,43
2002,43
2003,43
2004,43
2005,43
2006,43
2007,43
2008,43
2009,43
2010,43
2011,43
2012,43
2013,43
2014,43
2015,43
2016,43
2017,43
2018,43
2019,43
2020,43
2021,43
2022,43
2023,43
2024,44
2025,44
2026,44
2027,44
2028,44
2029,44
2030,44
2031,44
2032,44
2033,44
2034,44
2035,44
2036,44
2037,44
2038,44
2039,44
2040,44
2041,44
2042,44
2043,44
2044,44
2045,44
2046,44
2047,44
2048,44
2049,44
2050,44
2051,44
2052,44
2053,44
2054,44
2055,44
2056,44
2057,44
2058,44
2059,44
2060,44
2061,44
2062,44
2063,44
2064,44
2065,44
2066,44
2067,44
2068,44
2069,44
2070,45
2071,45
2072,45
2073,45
2074,45
2075,45
2076,45
2077,45
2078,45
2079,45
2080,45
2081,45
2082,45
2083,45
2084,45
2085,45
2086,45
2087,45
2088,45
2089,45
2090,45
2091,45
2092,45
2093,45
2094,45
2095,45
2096,45
2097,45
2098,45
2099,45
2100,45
2101,45
2102,45
2103,45
2104,45
2105,45
2106,45
2107,45
2108,45
2109,45
2110,45
2111,45
2112,45
2113,45
2114,45
2115,45
2116,46
2117,46
2118,46
2119,46
2120,46
2121,46
2122,46
2123,46
2124,46
2125,46
2126,46
2127,46
2128,46
2129,46
2130,46
2131,46
2132,46
2133,46
2134,46
2135,46
2136,46
2137,46
2138,46
2139,46
2140,46
2141,46
2142,46
2143,46
2144,46
2145,46
2146,46
2147,46
2148,46
2149,46
2150,46
2151,46
2152,46
2153,46
2154,46
2155,46
2156,46
2157,46
2158,46
2159,46
2160,46
2161,46
2162,47
2163,47
2164,47
2165,47
2166,47
2167,47
2168,47
2169,47
2170,47
2171,47
2172,47
2173,47
2174,47
2175,47
2176,47
2177,47
2178,47
2179,47
2180,47
2181,47
2182,47
2183,47
2184,47
2185,47
2186,47
2187,47
2188,47
2189,47
2190,47
2191,47
2192,47
2193,47
2194,47
2195,47
2196,47
2197,47
2198,47
2199,47
2200,47
2201,47
2202,47
2203,47
2204,47
2205,47
2206,47
2207,47
2208,48
2209,48
2210,48
2211,48
2212,48
2213,48
2214,48
2215,48
2216,48
2217,48
2218,48
2219,48
2220,48
2221,48
2222,48
2223,48
2224,48
2225,48
2226,48
2227,48
2228,48
2229,48
2230,48
2231,48
2232,48
2233,48
2234,48
2235,48
2236,48
2237,48
2238,48
2239,48
2240,48
2241,48
2242,48
2243,48
2244,48
2245,48
2246,48
2247,48
2248,48
2249,48
2250,48
2251,48
2252,48
2253,48
2254,49
2255,49
2256,49
2257,49
2258,49
2259,49
2260,49
2261,49
2262,49
2263,49
2264,49
2265,49
2266,49
2267,49
2268,49
2269,49
2270,49
2271,49
2272,49
2273,49
2274,49
2275,49
2276,49
2277,49
2278,49
2279,49
2280,49
2281,49
2282,49
2283,49
2284,49
2285,49
2286,49
2287,49
2288,49
2289,49
2290,49
2291,49
2292,49
2293,49
2294,49
2295,49
2296,49
2297,49
2298,49
2299,49
2300,50
2301,50
2302,50
2303,50
2304,50
2305,50
2306,50
2307,50
2308,50
2309,50
2310,50
2311,50
2312,50
2313,50
2314,50
2315,50
2316,50
2317,50
2318,50
2319,50
2320,50
2321,50
2322,50
2323,50
2324,50
2325,50
2326,50
2327,50
2328,50
2329,50
2330,50
2331,50
2332,50
2333,50
2334,50
2335,50
2336,50
2337,50
2338,50
2339,50
2340,50
2341,50
2342,50
2343,50
2344,50
2345,50
2346,51
2347,51
2348,51
2349,51
2350,51
2351,51
2352,51
2353,51
2354,51
2355,51
2356,51
2357,51
2358,51
2359,51
2360,51
2361,51
2362,51
2363,51
2364,51
2365,51
2366,51
2367,51
2368,51
2369,51
2370,51
2371,51
2372,51
2373,51
2374,51
2375,51
2376,51
2377,51
2378,51
2379,51
2380,51
2381,51
2382,51
2383,51
2384,51
2385,51
2386,51
2387,51
2388,51
2389,51
2390,51
2391,51
2392,52
2393,52
2394,52
2395,52
2396,52
2397,52
2398,52
2399,52
2400,52
2401,52
2402,52
2403,52
2404,52
2405,52
2406,52
2407,52
2408,52
2409,52
2410,52
2411,52
2412,52
2413,52
2414,52
2415,52
2416,52
2417,52
2418,52
2419,52
2420,52
2421,52
2422,52
2423,52
2424,52
2425,52
2426,52
2427,52
2428,52
2429,52
2430,52
2431,52
2432,52
2433,52
2434,52
2435,52
2436,52
2437,52
2438,53
2439,53
2440,53
2441,53
2442,53
2443,53
2444,53
2445,53
2446,53
2447,53
2448,53
2449,53
2450,53
2451,53
2452,53
2453,53
2454,53
2455,53
2456,53
2457,53
2458,53
2459,53
2460,53
2461,53
2462,53
2463,53
2464,53
2465,53
2466,53
2467,53
2468,53
2469,53
2470,53
2471,53
2472,53
2473,53
2474,53
2475,53
2476,53
2477,53
2478,53
2479,53
2480,53
2481,53
2482,53
2483,53
2484,54
2485,54
2486,54
2487,54
2488,54
2489,54
2490,54
2491,54
2492,54
2493,54
2494,54
2495,54
2496,54
2497,54
2498,54
2499,54
2500,54
2501,54
2502,54
2503,54
2504,54
2505,54
2506,54
2507,54
2508,54
2509,54
2510,54
2511,54
2512,54
2513,54
2514,54
2515,54
2516,54
2517,54
2518,54
2519,54
2520,54
2521,54
2522,54
2523,54
2524,54
2525,54
2526,54
2527,54
2528,54
2529,54
2530,55
2531,55
2532,55
2533,55
2534,55
2535,55
2536,55
2537,55
2538,55
2539,55
2540,55
2541,55
2542,55
2543,55
2544,55
2545,55
2546,55
2547,55
2548,55
2549,55
2550,55
2551,55
2552,55
2553,55
2554,55
2555,55
2556,55
2557,55
2558,55
2559,55
2560,55
2561,55
2562,55
2563,55
2564,55
2565,55
2566,55
2567,55
2568,55
2569,55
2570,55
2571,55
2572,55
2573,55
2574,55
2575,55
2576,56
2577,56
2578,56
2579,56
2580,56
2581,56
2582,56
2583,56
2584,56
2585,56
2586,56
2587,56
2588,56
2589,56
2590,56
2591,56
2592,56
2593,56
2594,56
2595,56
2596,56
2597,56
2598,56
2599,56
2600,56
2601,56
2602,56
2603,56
2604,56
2605,56
2606,56
2607,56
2608,56
2609,56
2610,56
2611,56
2612,56
2613,56
2614,56
2615,56
2616,56
2617,56
2618,56
2619,56
2620,56
2621,56
2622,57
2623,57
2624,57
2625,57
2626,57
2627,57
2628,57
2629,57
2630,57
2631,57
2632,57
2633,57
2634,57
2635,57
2636,57
2637,57
2638,57
2639,57
2640,57
2641,57
2642,57
2643,57
2644,57
2645,57
2646,57
2647,57
2648,57
2649,57
2650,57
2651,57
2652,57
2653,57
2654,57
2655,57
2656,57
2657,57
2658,57
2659,57
2660,57
2661,57
2662,57
2663,57
2664,57
2665,57
2666,57
2667,57
2668,58
2669,58
2670,58
2671,58
2672,58
2673,58
2674,58
2675,58
2676,58
2677,58
2678,58
2679,58
2680,58
2681,58
2682,58
2683,58
2684,58
2685,58
2686,58
2687,58
2688,58
2689,58
2690,58
2691,58
2692,58
2693,58
2694,58
2695,58
2696,58
2697,58
2698,58
2699,58
2700,58
2701,58
2702,58
2703,58
2704,58
2705,58
2706,58
2707,58
2708,58
2709,58
2710,58
2711,58
2712,58
2713,58
2714,59
2715,59
2716,59
2717,59
2718,59
2719,59
2720,59
2721,59
2722,59
2723,59
2724,59
2725,59
2726,59
2727,59
2728,59
2729,59
2730,59
2731,59
2732,59
2733,59
2734,59
2735,59
2736,59
2737,59
2738,59
2739,59
2740,59
2741,59
2742,59
2743,59
2744,59
2745,59
2746,59
2747,59
2748,59
2749,59
2750,59
2751,59
2752,59
2753,59
2754,59
2755,59
2756,59
2757,59
2758,59
2759,59
2760,60
2761,60
2762,60
2763,60
2764,60
2765,60
2766,60
2767,60
2768,60
2769,60
2770,60
2771,60
2772,60
2773,60
2774,60
2775,60
2776,60
2777,60
2778,60
2779,60
2780,60
2781,60
2782,60
2783,60
2784,60
2785,60
2786,60
2787,60
2788,60
2789,60
2790,60
2791,60
2792,60
2793,60
2794,60
2795,60
2796,60
2797,60
2798,60
2799,60
2800,60
2801,60
2802,60
2803,60
2804,60
2805,60
2806,61
2807,61
2808,61
2809,61
2810,61
2811,61
2812,61
2813,61
2814,61
2815,61
2816,61
2817,61
2818,61
2819,61
2820,61
2821,61
2822,61
2823,61
2824,61
2825,61
2826,61
2827,61
2828,61
2829,61
2830,61
2831,61
2832,61
2833,61
2834,61
2835,61
2836,61
2837,61
2838,61
2839,61
2840,61
2841,61
2842,61
2843,61
2844,61
2845,61
2846,61
2847,61
2848,61
2849,61
2850,61
2851,61
2852,62
2853,62
2854,62
2855,62
2856,62
2857,62
2858,62
2859,62
2860,62
2861,62
2862,62
2863,62
2864,62
2865,62
2866,62
2867,62
2868,62
2869,62
2870,62
2871,62
2872,62
2873,62
2874,62
2875,62
2876,62
2877,62
2878,62
2879,62
2880,62
2881,62
2882,62
2883,62
2884,62
2885,62
2886,62
2887,62
2888,62
2889,62
2890,62
2891,62
2892,62
2893,62
2894,62
2895,62
2896,62
2897,62
2898,63
2899,63
2900,63
2901,63
2902,63
2903,63
2904,63
2905,63
2906,63
2907,63
2908,63
2909,63
2910,63
2911,63
2912,63
2913,63
2914,63
2915,63
2916,63
2917,63
2918,63
2919,63
2920,63
2921,63
2922,63
2923,63
2924,63
2925,63
2926,63
2927,63
2928,63
2929,63
2930,63
2931,63
2932,63
2933,63
2934,63
2935,63
2936,63
2937,63
2938,63
2939,63
2940,63
2941,63
2942,63
2943,63
2944,64
2945,64
2946,64
2947,64
2948,64
2949,64
2950,64
2951,64
2952,64
2953,64
2954,64
2955,64
2956,64
2957,64
2958,64
2959,64
2960,64
2961,64
2962,64
2963,64
2964,64
2965,64
2966,64
2967,64
2968,64
2969,64
2970,64
2971,64
2972,64
2973,64
2974,64
2975,64
2976,64
2977,64
2978,64
2979,64
2980,64
2981,64
2982,64
2983,64
2984,64
2985,64
2986,64
2987,64
2988,64
2989,64
2990,65
2991,65
2992,65
2993,65
2994,65
2995,65
2996,65
2997,65
2998,65
2999,65
3000,65
3001,65
3002,65
3003,65
3004,65
3005,65
3006,65
3007,65
3008,65
3009,65
3010,65
3011,65
3012,65
3013,65
3014,65
3015,65
3016,65
3017,65
3018,65
3019,65
3020,65
3021,65
3022,65
3023,65
3024,65
3025,65
3026,65
3027,65
3028,65
3029,65
3030,65
3031,65
3032,65
3033,65
3034,65
3035,65
3036,66
3037,66
3038,66
3039,66
3040,66
3041,66
3042,66
3043,66
3044,66
3045,66
3046,66
3047,66
3048,66
3049,66
3050,66
3051,66
3052,66
3053,66
3054,66
3055,66
3056,66
3057,66
3058,66
3059,66
3060,66
3061,66
3062,66
3063,66
3064,66
3065,66
3066,66
3067,66
3068,66
3069,66
3070,66
3071,66
3072,66
3073,66
3074,66
3075,66
3076,66
3077,66
3078,66
3079,66
3080,66
3081,66
3082,67
3083,67
3084,67
3085,67
3086,67
3087,67
3088,67
3089,67
3090,67
3091,67
3092,67
3093,67
3094,67
3095,67
3096,67
3097,67
3098,67
3099,67
3100,67
3101,67
3102,67
3103,67
3104,67
3105,67
3106,67
3107,67
3108,67
3109,67
3110,67
3111,67
3112,67
3113,67
3114,67
3115,67
3116,67
3117,67
3118,67
3119,67
3120,67
3121,67
3122,67
3123,67
3124,67
3125,67
3126,67
3127,67
