0,0
1,0
2,0
3,0
4,0
5,0
6,0
7,0
8,0
9,0
10,0
11,0
12,0
13,0
14,0
15,0
16,0
17,0
18,0
19,0
20,0
21,0
22,0
23,0
24,0
25,0
26,0
27,0
28,1
29,1
30,1
31,1
32,1
33,1
34,1
35,1
36,1
37,1
38,1
39,1
40,1
41,1
42,1
43,1
44,1
45,1
46,1
47,1
48,1
49,1
50,1
51,1
52,1
53,1
54,1
55,1
56,2
57,2
58,2
59,2
60,2
61,2
62,2
63,2
64,2
65,2
66,2
67,2
68,2
69,2
70,2
71,2
72,2
73,2
74,2
75,2
76,2
77,2
78,2
79,2
80,2
81,2
82,2
83,2
84,3
85,3
86,3
87,3
88,3
89,3
90,3
91,3
92,3
93,3
94,3
95,3
96,3
97,3
98,3
99,3
100,3
101,3
102,3
103,3
104,3
105,3
106,3
107,3
108,3
109,3
110,3
111,3
112,4
113,4
114,4
115,4
116,4
117,4
118,4
119,4
120,4
121,4
122,4
123,4
124,4
125,4
126,4
127,4
128,4
129,4
130,4
131,4
132,4
133,4
134,4
135,4
136,4
137,4
138,4
139,4
140,5
141,5
142,5
143,5
144,5
145,5
146,5
147,5
148,5
149,5
150,5
151,5
152,5
153,5
154,5
155,5
156,5
157,5
158,5
159,5
160,5
161,5
162,5
163,5
164,5
165,5
166,5
167,5
168,6
169,6
170,6
171,6
172,6
173,6
174,6
175,6
176,6
177,6
178,6
179,6
180,6
181,6
182,6
183,6
184,6
185,6
186,6
187,6
188,6
189,6
190,6
191,6
192,6
193,6
194,6
195,6
196,7
197,7
198,7
199,7
200,7
201,7
202,7
203,7
204,7
205,7
206,7
207,7
208,7
209,7
210,7
211,7
212,7
213,7
214,7
215,7
216,7
217,7
218,7
219,7
220,7
221,7
222,7
223,7
224,8
225,8
226,8
227,8
228,8
229,8
230,8
231,8
232,8
233,8
234,8
235,8
236,8
237,8
238,8
239,8
240,8
241,8
242,8
243,8
244,8
245,8
246,8
247,8
248,8
249,8
250,8
251,8
252,9
253,9
254,9
255,9
256,9
257,9
258,9
259,9
260,9
261,9
262,9
263,9
264,9
265,9
266,9
267,9
268,9
269,9
270,9
271,9
272,9
273,9
274,9
275,9
276,9
277,9
278,9
279,9
280,10
281,10
282,10
283,10
284,10
285,10
286,10
287,10
288,10
289,10
290,10
291,10
292,10
293,10
294,10
295,10
296,10
297,10
298,10
299,10
300,10
301,10
302,10
303,10
304,10
305,10
306,10
307,10
308,11
309,11
310,11
311,11
312,11
313,11
314,11
315,11
316,11
317,11
318,11
319,11
320,11
321,11
322,11
323,11
324,11
325,11
326,11
327,11
328,11
329,11
330,11
331,11
332,11
333,11
334,11
335,11
336,12
337,12
338,12
339,12
340,12
341,12
342,12
343,12
344,12
345,12
346,12
347,12
348,12
349,12
350,12
351,12
352,12
353,12
354,12
355,12
356,12
357,12
358,12
359,12
360,12
361,12
362,12
363,12
364,12
365,13
366,13
367,13
368,13
369,13
370,13
371,13
372,13
373,13
374,13
375,13
376,13
377,13
378,13
379,13
380,13
381,13
382,13
383,13
384,13
385,13
386,13
387,13
388,13
389,13
390,13
391,13
392,13
393,13
394,14
395,14
396,14
397,14
398,14
399,14
400,14
401,14
402,14
403,14
404,14
405,14
406,14
407,14
408,14
409,14
410,14
411,14
412,14
413,14
414,14
415,14
416,14
417,14
418,14
419,14
420,14
421,14
422,14
423,15
424,15
425,15
426,15
427,15
428,15
429,15
430,15
431,15
432,15
433,15
434,15
435,15
436,15
437,15
438,15
439,15
440,15
441,15
442,15
443,15
444,15
445,15
446,15
447,15
448,15
449,15
450,15
451,15
452,16
453,16
454,16
455,16
456,16
457,16
458,16
459,16
460,16
461,16
462,16
463,16
464,16
465,16
466,16
467,16
468,16
469,16
470,16
471,16
472,16
473,16
474,16
475,16
476,16
477,16
478,16
479,16
480,16
481,17
482,17
483,17
484,17
485,17
486,17
487,17
488,17
489,17
490,17
491,17
492,17
493,17
494,17
495,17
496,17
497,17
498,17
499,17
500,17
501,17
502,17
503,17
504,17
505,17
506,17
507,17
508,17
509,17
510,18
511,18
512,18
513,18
514,18
515,18
516,18
517,18
518,18
519,18
520,18
521,18
522,18
523,18
524,18
525,18
526,18
527,18
528,18
529,18
530,18
531,18
532,18
533,18
534,18
535,18
536,18
537,18
538,18
539,19
540,19
541,19
542,19
543,19
544,19
545,19
546,19
547,19
548,19
549,19
550,19
551,19
552,19
553,19
554,19
555,19
556,19
557,19
558,19
559,19
560,19
561,19
562,19
563,19
564,19
565,19
566,19
567,19
568,20
569,20
570,20
571,20
572,20
573,20
574,20
575,20
576,20
577,20
578,20
579,20
580,20
581,20
582,20
583,20
584,20
585,20
586,20
587,20
588,20
589,20
590,20
591,20
592,20
593,20
594,20
595,20
596,20
597,21
598,21
599,21
600,21
601,21
602,21
603,21
604,21
605,21
606,21
607,21
608,21
609,21
610,21
611,21
612,21
613,21
614,21
615,21
616,21
617,21
618,21
619,21
620,21
621,21
622,21
623,21
624,21
625,21
626,22
627,22
628,22
629,22
630,22
631,22
632,22
633,22
634,22
635,22
636,22
637,22
638,22
639,22
640,22
641,22
642,22
643,22
644,22
645,22
646,22
647,22
648,22
649,22
650,22
651,22
652,22
653,22
654,22
655,23
656,23
657,23
658,23
659,23
660,23
661,23
662,23
663,23
664,23
665,23
666,23
667,23
668,23
669,23
670,23
671,23
672,23
673,23
674,23
675,23
676,23
677,23
678,23
679,23
680,23
681,23
682,23
683,23
684,24
685,24
686,24
687,24
688,24
689,24
690,24
691,24
692,24
693,24
694,24
695,24
696,24
697,24
698,24
699,24
700,24
701,24
702,24
703,24
704,24
705,24
706,24
707,24
708,24
709,24
710,24
711,24
712,24
713,25
714,25
715,25
716,25
717,25
718,25
719,25
720,25
721,25
722,25
723,25
724,25
725,25
726,25
727,25
728,25
729,25
730,25
731,25
732,25
733,25
734,25
735,25
736,25
737,25
738,25
739,25
740,25
741,25
742,26
743,26
744,26
745,26
746,26
747,26
748,26
749,26
750,26
751,26
752,26
753,26
754,26
755,26
756,26
757,26
758,26
759,26
760,26
761,26
762,26
763,26
764,26
765,26
766,26
767,26
768,26
769,26
770,26
771,27
772,27
773,27
774,27
775,27
776,27
777,27
778,27
779,27
780,27
781,27
782,27
783,27
784,27
785,27
786,27
787,27
788,27
789,27
790,27
791,27
792,27
793,27
794,27
795,27
796,27
797,27
798,27
799,27
800,28
801,28
802,28
803,28
804,28
805,28
806,28
807,28
808,28
809,28
810,28
811,28
812,28
813,28
814,28
815,28
816,28
817,28
818,28
819,28
820,28
821,28
822,28
823,28
824,28
825,28
826,28
827,28
828,28
829,29
830,29
831,29
832,29
833,29
834,29
835,29
836,29
837,29
838,29
839,29
840,29
841,29
842,29
843,29
844,29
845,29
846,29
847,29
848,29
849,29
850,29
851,29
852,29
853,29
854,29
855,29
856,29
857,29
858,30
859,30
860,30
861,30
862,30
863,30
864,30
865,30
866,30
867,30
868,30
869,30
870,30
871,30
872,30
873,30
874,30
875,30
876,30
877,30
878,30
879,30
880,30
881,30
882,30
883,30
884,30
885,30
886,30
887,31
888,31
889,31
890,31
891,31
892,31
893,31
894,31
895,31
896,31
897,31
898,31
899,31
900,31
901,31
902,31
903,31
904,31
905,31
906,31
907,31
908,31
909,31
910,31
911,31
912,31
913,31
914,31
915,31
916,32
917,32
918,32
919,32
920,32
921,32
922,32
923,32
924,32
925,32
926,32
927,32
928,32
929,32
930,32
931,32
932,32
933,32
934,32
935,32
936,32
937,32
938,32
939,32
940,32
941,32
942,32
943,32
944,32
945,33
946,33
947,33
948,33
949,33
950,33
951,33
952,33
953,33
954,33
955,33
956,33
957,33
958,33
959,33
960,33
961,33
962,33
963,33
964,33
965,33
966,33
967,33
968,33
969,33
970,33
971,33
972,33
973,33
974,34
975,34
976,34
977,34
978,34
979,34
980,34
981,34
982,34
983,34
984,34
985,34
986,34
987,34
988,34
989,34
990,34
991,34
992,34
993,34
994,34
995,34
996,34
997,34
998,34
999,34
1000,34
1001,34
1002,34
1003,35
1004,35
1005,35
1006,35
1007,35
1008,35
1009,35
1010,35
1011,35
1012,35
1013,35
1014,35
1015,35
1016,35
1017,35
1018,35
1019,35
1020,35
1021,35
1022,35
1023,35
1024,35
1025,35
1026,35
1027,35
1028,35
1029,35
1030,35
1031,35
1032,36
1033,36
1034,36
1035,36
1036,36
1037,36
1038,36
1039,36
1040,36
1041,36
1042,36
1043,36
1044,36
1045,36
1046,36
1047,36
1048,36
1049,36
1050,36
1051,36
1052,36
1053,36
1054,36
1055,36
1056,36
1057,36
1058,36
1059,36
1060,36
1061,37
1062,37
1063,37
1064,37
1065,37
1066,37
1067,37
1068,37
1069,37
1070,37
1071,37
1072,37
1073,37
1074,37
1075,37
1076,37
1077,37
1078,37
1079,37
1080,37
1081,37
1082,37
1083,37
1084,37
1085,37
1086,37
1087,37
1088,37
1089,37
1090,38
1091,38
1092,38
1093,38
1094,38
1095,38
1096,38
1097,38
1098,38
1099,38
1100,38
1101,38
1102,38
1103,38
1104,38
1105,38
1106,38
1107,38
1108,38
1109,38
1110,38
1111,38
1112,38
1113,38
1114,38
1115,38
1116,38
1117,38
1118,38
1119,39
1120,39
1121,39
1122,39
1123,39
1124,39
1125,39
1126,39
1127,39
1128,39
1129,39
1130,39
1131,39
1132,39
1133,39
1134,39
1135,39
1136,39
1137,39
1138,39
1139,39
1140,39
1141,39
1142,39
1143,39
1144,39
1145,39
1146,39
1147,39
1148,40
1149,40
1150,40
1151,40
1152,40
1153,40
1154,40
1155,40
1156,40
1157,40
1158,40
1159,40
1160,40
1161,40
1162,40
1163,40
1164,40
1165,40
1166,40
1167,40
1168,40
1169,40
1170,40
1171,40
1172,40
1173,40
1174,40
1175,40
1176,40
1177,41
1178,41
1179,41
1180,41
1181,41
1182,41
1183,41
1184,41
1185,41
1186,41
1187,41
1188,41
1189,41
1190,41
1191,41
1192,41
1193,41
1194,41
1195,41
1196,41
1197,41
1198,41
1199,41
1200,41
1201,41
1202,41
1203,41
1204,41
1205,41
1206,42
1207,42
1208,42
1209,42
1210,42
1211,42
1212,42
1213,42
1214,42
1215,42
1216,42
1217,42
1218,42
1219,42
1220,42
1221,42
1222,42
1223,42
1224,42
1225,42
1226,42
1227,42
1228,42
1229,42
1230,42
1231,42
1232,42
1233,42
1234,42
1235,43
1236,43
1237,43
1238,43
1239,43
1240,43
1241,43
1242,43
1243,43
1244,43
1245,43
1246,43
1247,43
1248,43
1249,43
1250,43
1251,43
1252,43
1253,43
1254,43
1255,43
1256,43
1257,43
1258,43
1259,43
1260,43
1261,43
1262,43
1263,43
1264,44
1265,44
1266,44
1267,44
1268,44
1269,44
1270,44
1271,44
1272,44
1273,44
1274,44
1275,44
1276,44
1277,44
1278,44
1279,44
1280,44
1281,44
1282,44
1283,44
1284,44
1285,44
1286,44
1287,44
1288,44
1289,44
1290,44
1291,44
1292,44
1293,45
1294,45
1295,45
1296,45
1297,45
1298,45
1299,45
1300,45
1301,45
1302,45
1303,45
1304,45
1305,45
1306,45
1307,45
1308,45
1309,45
1310,45
1311,45
1312,45
1313,45
1314,45
1315,45
1316,45
1317,45
1318,45
1319,45
1320,45
1321,45
1322,46
1323,46
1324,46
1325,46
1326,46
1327,46
1328,46
1329,46
1330,46
1331,46
1332,46
1333,46
1334,46
1335,46
1336,46
1337,46
1338,46
1339,46
1340,46
1341,46
1342,46
1343,46
1344,46
1345,46
1346,46
1347,46
1348,46
1349,46
1350,46
1351,47
1352,47
1353,47
1354,47
1355,47
1356,47
1357,47
1358,47
1359,47
1360,47
1361,47
1362,47
1363,47
1364,47
1365,47
1366,47
1367,47
1368,47
1369,47
1370,47
1371,47
1372,47
1373,47
1374,47
1375,47
1376,47
1377,47
1378,47
1379,47
1380,48
1381,48
1382,48
1383,48
1384,48
1385,48
1386,48
1387,48
1388,48
1389,48
1390,48
1391,48
1392,48
1393,48
1394,48
1395,48
1396,48
1397,48
1398,48
1399,48
1400,48
1401,48
1402,48
1403,48
1404,48
1405,48
1406,48
1407,48
1408,48
1409,49
1410,49
1411,49
1412,49
1413,49
1414,49
1415,49
1416,49
1417,49
1418,49
1419,49
1420,49
1421,49
1422,49
1423,49
1424,49
1425,49
1426,49
1427,49
1428,49
1429,49
1430,49
1431,49
1432,49
1433,49
1434,49
1435,49
1436,49
1437,49
1438,50
1439,50
1440,50
1441,50
1442,50
1443,50
1444,50
1445,50
1446,50
1447,50
1448,50
1449,50
1450,50
1451,50
1452,50
1453,50
1454,50
1455,50
1456,50
1457,50
1458,50
1459,50
1460,50
1461,50
1462,50
1463,50
1464,50
1465,50
1466,50
1467,51
1468,51
1469,51
1470,51
1471,51
1472,51
1473,51
1474,51
1475,51
1476,51
1477,51
1478,51
1479,51
1480,51
1481,51
1482,51
1483,51
1484,51
1485,51
1486,51
1487,51
1488,51
1489,51
1490,51
1491,51
1492,51
1493,51
1494,51
1495,51
1496,52
1497,52
1498,52
1499,52
1500,52
1501,52
1502,52
1503,52
1504,52
1505,52
1506,52
1507,52
1508,52
1509,52
1510,52
1511,52
1512,52
1513,52
1514,52
1515,52
1516,52
1517,52
1518,52
1519,52
1520,52
1521,52
1522,52
1523,52
1524,52
1525,53
1526,53
1527,53
1528,53
1529,53
1530,53
1531,53
1532,53
1533,53
1534,53
1535,53
1536,53
1537,53
1538,53
1539,53
1540,53
1541,53
1542,53
1543,53
1544,53
1545,53
1546,53
1547,53
1548,53
1549,53
1550,53
1551,53
1552,53
1553,53
1554,54
1555,54
1556,54
1557,54
1558,54
1559,54
1560,54
1561,54
1562,54
1563,54
1564,54
1565,54
1566,54
1567,54
1568,54
1569,54
1570,54
1571,54
1572,54
1573,54
1574,54
1575,54
1576,54
1577,54
1578,54
1579,54
1580,54
1581,54
1582,54
1583,55
1584,55
1585,55
1586,55
1587,55
1588,55
1589,55
1590,55
1591,55
1592,55
1593,55
1594,55
1595,55
1596,55
1597,55
1598,55
1599,55
1600,55
1601,55
1602,55
1603,55
1604,55
1605,55
1606,55
1607,55
1608,55
1609,55
1610,55
1611,55
1612,56
1613,56
1614,56
1615,56
1616,56
1617,56
1618,56
1619,56
1620,56
1621,56
1622,56
1623,56
1624,56
1625,56
1626,56
1627,56
1628,56
1629,56
1630,56
1631,56
1632,56
1633,56
1634,56
1635,56
1636,56
1637,56
1638,56
1639,56
1640,56
1641,57
1642,57
1643,57
1644,57
1645,57
1646,57
1647,57
1648,57
1649,57
1650,57
1651,57
1652,57
1653,57
1654,57
1655,57
1656,57
1657,57
1658,57
1659,57
1660,57
1661,57
1662,57
1663,57
1664,57
1665,57
1666,57
1667,57
1668,57
1669,57
1670,58
1671,58
1672,58
1673,58
1674,58
1675,58
1676,58
1677,58
1678,58
1679,58
1680,58
1681,58
1682,58
1683,58
1684,58
1685,58
1686,58
1687,58
1688,58
1689,58
1690,58
1691,58
1692,58
1693,58
1694,58
1695,58
1696,58
1697,58
1698,58
1699,59
1700,59
1701,59
1702,59
1703,59
1704,59
1705,59
1706,59
1707,59
1708,59
1709,59
1710,59
1711,59
1712,59
1713,59
1714,59
1715,59
1716,59
1717,59
1718,59
1719,59
1720,59
1721,59
1722,59
1723,59
1724,59
1725,59
1726,59
1727,59
