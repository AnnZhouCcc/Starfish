0,0
1,0
2,0
3,0
4,0
5,0
6,0
7,0
8,0
9,0
10,0
11,0
12,0
13,0
14,0
15,0
16,0
17,0
18,0
19,0
20,0
21,0
22,0
23,0
24,0
25,0
26,0
27,0
28,0
29,0
30,0
31,0
32,0
33,0
34,0
35,0
36,0
37,0
38,0
39,0
40,0
41,0
42,0
43,0
44,0
45,0
46,0
47,0
48,0
49,0
50,0
51,0
52,0
53,0
54,0
55,0
56,0
57,1
58,1
59,1
60,1
61,1
62,1
63,1
64,1
65,1
66,1
67,1
68,1
69,1
70,1
71,1
72,1
73,1
74,1
75,1
76,1
77,1
78,1
79,1
80,1
81,1
82,1
83,1
84,1
85,1
86,1
87,1
88,1
89,1
90,1
91,1
92,1
93,1
94,1
95,1
96,1
97,1
98,1
99,1
100,1
101,1
102,1
103,1
104,1
105,1
106,1
107,1
108,1
109,1
110,1
111,1
112,1
113,1
114,2
115,2
116,2
117,2
118,2
119,2
120,2
121,2
122,2
123,2
124,2
125,2
126,2
127,2
128,2
129,2
130,2
131,2
132,2
133,2
134,2
135,2
136,2
137,2
138,2
139,2
140,2
141,2
142,2
143,2
144,2
145,2
146,2
147,2
148,2
149,2
150,2
151,2
152,2
153,2
154,2
155,2
156,2
157,2
158,2
159,2
160,2
161,2
162,2
163,2
164,2
165,2
166,2
167,2
168,2
169,2
170,2
171,3
172,3
173,3
174,3
175,3
176,3
177,3
178,3
179,3
180,3
181,3
182,3
183,3
184,3
185,3
186,3
187,3
188,3
189,3
190,3
191,3
192,3
193,3
194,3
195,3
196,3
197,3
198,3
199,3
200,3
201,3
202,3
203,3
204,3
205,3
206,3
207,3
208,3
209,3
210,3
211,3
212,3
213,3
214,3
215,3
216,3
217,3
218,3
219,3
220,3
221,3
222,3
223,3
224,3
225,3
226,3
227,3
228,4
229,4
230,4
231,4
232,4
233,4
234,4
235,4
236,4
237,4
238,4
239,4
240,4
241,4
242,4
243,4
244,4
245,4
246,4
247,4
248,4
249,4
250,4
251,4
252,4
253,4
254,4
255,4
256,4
257,4
258,4
259,4
260,4
261,4
262,4
263,4
264,4
265,4
266,4
267,4
268,4
269,4
270,4
271,4
272,4
273,4
274,4
275,4
276,4
277,4
278,4
279,4
280,4
281,4
282,4
283,4
284,4
285,5
286,5
287,5
288,5
289,5
290,5
291,5
292,5
293,5
294,5
295,5
296,5
297,5
298,5
299,5
300,5
301,5
302,5
303,5
304,5
305,5
306,5
307,5
308,5
309,5
310,5
311,5
312,5
313,5
314,5
315,5
316,5
317,5
318,5
319,5
320,5
321,5
322,5
323,5
324,5
325,5
326,5
327,5
328,5
329,5
330,5
331,5
332,5
333,5
334,5
335,5
336,5
337,5
338,5
339,5
340,5
341,5
342,6
343,6
344,6
345,6
346,6
347,6
348,6
349,6
350,6
351,6
352,6
353,6
354,6
355,6
356,6
357,6
358,6
359,6
360,6
361,6
362,6
363,6
364,6
365,6
366,6
367,6
368,6
369,6
370,6
371,6
372,6
373,6
374,6
375,6
376,6
377,6
378,6
379,6
380,6
381,6
382,6
383,6
384,6
385,6
386,6
387,6
388,6
389,6
390,6
391,6
392,6
393,6
394,6
395,6
396,6
397,6
398,6
399,7
400,7
401,7
402,7
403,7
404,7
405,7
406,7
407,7
408,7
409,7
410,7
411,7
412,7
413,7
414,7
415,7
416,7
417,7
418,7
419,7
420,7
421,7
422,7
423,7
424,7
425,7
426,7
427,7
428,7
429,7
430,7
431,7
432,7
433,7
434,7
435,7
436,7
437,7
438,7
439,7
440,7
441,7
442,7
443,7
444,7
445,7
446,7
447,7
448,7
449,7
450,7
451,7
452,7
453,7
454,7
455,7
456,8
457,8
458,8
459,8
460,8
461,8
462,8
463,8
464,8
465,8
466,8
467,8
468,8
469,8
470,8
471,8
472,8
473,8
474,8
475,8
476,8
477,8
478,8
479,8
480,8
481,8
482,8
483,8
484,8
485,8
486,8
487,8
488,8
489,8
490,8
491,8
492,8
493,8
494,8
495,8
496,8
497,8
498,8
499,8
500,8
501,8
502,8
503,8
504,8
505,8
506,8
507,8
508,8
509,8
510,8
511,8
512,8
513,9
514,9
515,9
516,9
517,9
518,9
519,9
520,9
521,9
522,9
523,9
524,9
525,9
526,9
527,9
528,9
529,9
530,9
531,9
532,9
533,9
534,9
535,9
536,9
537,9
538,9
539,9
540,9
541,9
542,9
543,9
544,9
545,9
546,9
547,9
548,9
549,9
550,9
551,9
552,9
553,9
554,9
555,9
556,9
557,9
558,9
559,9
560,9
561,9
562,9
563,9
564,9
565,9
566,9
567,9
568,9
569,9
570,10
571,10
572,10
573,10
574,10
575,10
576,10
577,10
578,10
579,10
580,10
581,10
582,10
583,10
584,10
585,10
586,10
587,10
588,10
589,10
590,10
591,10
592,10
593,10
594,10
595,10
596,10
597,10
598,10
599,10
600,10
601,10
602,10
603,10
604,10
605,10
606,10
607,10
608,10
609,10
610,10
611,10
612,10
613,10
614,10
615,10
616,10
617,10
618,10
619,10
620,10
621,10
622,10
623,10
624,10
625,10
626,10
627,11
628,11
629,11
630,11
631,11
632,11
633,11
634,11
635,11
636,11
637,11
638,11
639,11
640,11
641,11
642,11
643,11
644,11
645,11
646,11
647,11
648,11
649,11
650,11
651,11
652,11
653,11
654,11
655,11
656,11
657,11
658,11
659,11
660,11
661,11
662,11
663,11
664,11
665,11
666,11
667,11
668,11
669,11
670,11
671,11
672,11
673,11
674,11
675,11
676,11
677,11
678,11
679,11
680,11
681,11
682,11
683,11
684,12
685,12
686,12
687,12
688,12
689,12
690,12
691,12
692,12
693,12
694,12
695,12
696,12
697,12
698,12
699,12
700,12
701,12
702,12
703,12
704,12
705,12
706,12
707,12
708,12
709,12
710,12
711,12
712,12
713,12
714,12
715,12
716,12
717,12
718,12
719,12
720,12
721,12
722,12
723,12
724,12
725,12
726,12
727,12
728,12
729,12
730,12
731,12
732,12
733,12
734,12
735,12
736,12
737,12
738,12
739,12
740,12
741,13
742,13
743,13
744,13
745,13
746,13
747,13
748,13
749,13
750,13
751,13
752,13
753,13
754,13
755,13
756,13
757,13
758,13
759,13
760,13
761,13
762,13
763,13
764,13
765,13
766,13
767,13
768,13
769,13
770,13
771,13
772,13
773,13
774,13
775,13
776,13
777,13
778,13
779,13
780,13
781,13
782,13
783,13
784,13
785,13
786,13
787,13
788,13
789,13
790,13
791,13
792,13
793,13
794,13
795,13
796,13
797,13
798,14
799,14
800,14
801,14
802,14
803,14
804,14
805,14
806,14
807,14
808,14
809,14
810,14
811,14
812,14
813,14
814,14
815,14
816,14
817,14
818,14
819,14
820,14
821,14
822,14
823,14
824,14
825,14
826,14
827,14
828,14
829,14
830,14
831,14
832,14
833,14
834,14
835,14
836,14
837,14
838,14
839,14
840,14
841,14
842,14
843,14
844,14
845,14
846,14
847,14
848,14
849,14
850,14
851,14
852,14
853,14
854,14
855,15
856,15
857,15
858,15
859,15
860,15
861,15
862,15
863,15
864,15
865,15
866,15
867,15
868,15
869,15
870,15
871,15
872,15
873,15
874,15
875,15
876,15
877,15
878,15
879,15
880,15
881,15
882,15
883,15
884,15
885,15
886,15
887,15
888,15
889,15
890,15
891,15
892,15
893,15
894,15
895,15
896,15
897,15
898,15
899,15
900,15
901,15
902,15
903,15
904,15
905,15
906,15
907,15
908,15
909,15
910,15
911,15
912,16
913,16
914,16
915,16
916,16
917,16
918,16
919,16
920,16
921,16
922,16
923,16
924,16
925,16
926,16
927,16
928,16
929,16
930,16
931,16
932,16
933,16
934,16
935,16
936,16
937,16
938,16
939,16
940,16
941,16
942,16
943,16
944,16
945,16
946,16
947,16
948,16
949,16
950,16
951,16
952,16
953,16
954,16
955,16
956,16
957,16
958,16
959,16
960,16
961,16
962,16
963,16
964,16
965,16
966,16
967,16
968,16
969,17
970,17
971,17
972,17
973,17
974,17
975,17
976,17
977,17
978,17
979,17
980,17
981,17
982,17
983,17
984,17
985,17
986,17
987,17
988,17
989,17
990,17
991,17
992,17
993,17
994,17
995,17
996,17
997,17
998,17
999,17
1000,17
1001,17
1002,17
1003,17
1004,17
1005,17
1006,17
1007,17
1008,17
1009,17
1010,17
1011,17
1012,17
1013,17
1014,17
1015,17
1016,17
1017,17
1018,17
1019,17
1020,17
1021,17
1022,17
1023,17
1024,17
1025,17
1026,18
1027,18
1028,18
1029,18
1030,18
1031,18
1032,18
1033,18
1034,18
1035,18
1036,18
1037,18
1038,18
1039,18
1040,18
1041,18
1042,18
1043,18
1044,18
1045,18
1046,18
1047,18
1048,18
1049,18
1050,18
1051,18
1052,18
1053,18
1054,18
1055,18
1056,18
1057,18
1058,18
1059,18
1060,18
1061,18
1062,18
1063,18
1064,18
1065,18
1066,18
1067,18
1068,18
1069,18
1070,18
1071,18
1072,18
1073,18
1074,18
1075,18
1076,18
1077,18
1078,18
1079,18
1080,18
1081,18
1082,18
1083,19
1084,19
1085,19
1086,19
1087,19
1088,19
1089,19
1090,19
1091,19
1092,19
1093,19
1094,19
1095,19
1096,19
1097,19
1098,19
1099,19
1100,19
1101,19
1102,19
1103,19
1104,19
1105,19
1106,19
1107,19
1108,19
1109,19
1110,19
1111,19
1112,19
1113,19
1114,19
1115,19
1116,19
1117,19
1118,19
1119,19
1120,19
1121,19
1122,19
1123,19
1124,19
1125,19
1126,19
1127,19
1128,19
1129,19
1130,19
1131,19
1132,19
1133,19
1134,19
1135,19
1136,19
1137,19
1138,19
1139,19
1140,20
1141,20
1142,20
1143,20
1144,20
1145,20
1146,20
1147,20
1148,20
1149,20
1150,20
1151,20
1152,20
1153,20
1154,20
1155,20
1156,20
1157,20
1158,20
1159,20
1160,20
1161,20
1162,20
1163,20
1164,20
1165,20
1166,20
1167,20
1168,20
1169,20
1170,20
1171,20
1172,20
1173,20
1174,20
1175,20
1176,20
1177,20
1178,20
1179,20
1180,20
1181,20
1182,20
1183,20
1184,20
1185,20
1186,20
1187,20
1188,20
1189,20
1190,20
1191,20
1192,20
1193,20
1194,20
1195,20
1196,20
1197,21
1198,21
1199,21
1200,21
1201,21
1202,21
1203,21
1204,21
1205,21
1206,21
1207,21
1208,21
1209,21
1210,21
1211,21
1212,21
1213,21
1214,21
1215,21
1216,21
1217,21
1218,21
1219,21
1220,21
1221,21
1222,21
1223,21
1224,21
1225,21
1226,21
1227,21
1228,21
1229,21
1230,21
1231,21
1232,21
1233,21
1234,21
1235,21
1236,21
1237,21
1238,21
1239,21
1240,21
1241,21
1242,21
1243,21
1244,21
1245,21
1246,21
1247,21
1248,21
1249,21
1250,21
1251,21
1252,21
1253,21
1254,22
1255,22
1256,22
1257,22
1258,22
1259,22
1260,22
1261,22
1262,22
1263,22
1264,22
1265,22
1266,22
1267,22
1268,22
1269,22
1270,22
1271,22
1272,22
1273,22
1274,22
1275,22
1276,22
1277,22
1278,22
1279,22
1280,22
1281,22
1282,22
1283,22
1284,22
1285,22
1286,22
1287,22
1288,22
1289,22
1290,22
1291,22
1292,22
1293,22
1294,22
1295,22
1296,22
1297,22
1298,22
1299,22
1300,22
1301,22
1302,22
1303,22
1304,22
1305,22
1306,22
1307,22
1308,22
1309,22
1310,22
1311,23
1312,23
1313,23
1314,23
1315,23
1316,23
1317,23
1318,23
1319,23
1320,23
1321,23
1322,23
1323,23
1324,23
1325,23
1326,23
1327,23
1328,23
1329,23
1330,23
1331,23
1332,23
1333,23
1334,23
1335,23
1336,23
1337,23
1338,23
1339,23
1340,23
1341,23
1342,23
1343,23
1344,23
1345,23
1346,23
1347,23
1348,23
1349,23
1350,23
1351,23
1352,23
1353,23
1354,23
1355,23
1356,23
1357,23
1358,23
1359,23
1360,23
1361,23
1362,23
1363,23
1364,23
1365,23
1366,23
1367,23
1368,24
1369,24
1370,24
1371,24
1372,24
1373,24
1374,24
1375,24
1376,24
1377,24
1378,24
1379,24
1380,24
1381,24
1382,24
1383,24
1384,24
1385,24
1386,24
1387,24
1388,24
1389,24
1390,24
1391,24
1392,24
1393,24
1394,24
1395,24
1396,24
1397,24
1398,24
1399,24
1400,24
1401,24
1402,24
1403,24
1404,24
1405,24
1406,24
1407,24
1408,24
1409,24
1410,24
1411,24
1412,24
1413,24
1414,24
1415,24
1416,24
1417,24
1418,24
1419,24
1420,24
1421,24
1422,24
1423,24
1424,24
1425,25
1426,25
1427,25
1428,25
1429,25
1430,25
1431,25
1432,25
1433,25
1434,25
1435,25
1436,25
1437,25
1438,25
1439,25
1440,25
1441,25
1442,25
1443,25
1444,25
1445,25
1446,25
1447,25
1448,25
1449,25
1450,25
1451,25
1452,25
1453,25
1454,25
1455,25
1456,25
1457,25
1458,25
1459,25
1460,25
1461,25
1462,25
1463,25
1464,25
1465,25
1466,25
1467,25
1468,25
1469,25
1470,25
1471,25
1472,25
1473,25
1474,25
1475,25
1476,25
1477,25
1478,25
1479,25
1480,25
1481,25
1482,26
1483,26
1484,26
1485,26
1486,26
1487,26
1488,26
1489,26
1490,26
1491,26
1492,26
1493,26
1494,26
1495,26
1496,26
1497,26
1498,26
1499,26
1500,26
1501,26
1502,26
1503,26
1504,26
1505,26
1506,26
1507,26
1508,26
1509,26
1510,26
1511,26
1512,26
1513,26
1514,26
1515,26
1516,26
1517,26
1518,26
1519,26
1520,26
1521,26
1522,26
1523,26
1524,26
1525,26
1526,26
1527,26
1528,26
1529,26
1530,26
1531,26
1532,26
1533,26
1534,26
1535,26
1536,26
1537,26
1538,26
1539,27
1540,27
1541,27
1542,27
1543,27
1544,27
1545,27
1546,27
1547,27
1548,27
1549,27
1550,27
1551,27
1552,27
1553,27
1554,27
1555,27
1556,27
1557,27
1558,27
1559,27
1560,27
1561,27
1562,27
1563,27
1564,27
1565,27
1566,27
1567,27
1568,27
1569,27
1570,27
1571,27
1572,27
1573,27
1574,27
1575,27
1576,27
1577,27
1578,27
1579,27
1580,27
1581,27
1582,27
1583,27
1584,27
1585,27
1586,27
1587,27
1588,27
1589,27
1590,27
1591,27
1592,27
1593,27
1594,27
1595,27
1596,28
1597,28
1598,28
1599,28
1600,28
1601,28
1602,28
1603,28
1604,28
1605,28
1606,28
1607,28
1608,28
1609,28
1610,28
1611,28
1612,28
1613,28
1614,28
1615,28
1616,28
1617,28
1618,28
1619,28
1620,28
1621,28
1622,28
1623,28
1624,28
1625,28
1626,28
1627,28
1628,28
1629,28
1630,28
1631,28
1632,28
1633,28
1634,28
1635,28
1636,28
1637,28
1638,28
1639,28
1640,28
1641,28
1642,28
1643,28
1644,28
1645,28
1646,28
1647,28
1648,28
1649,28
1650,28
1651,28
1652,28
1653,29
1654,29
1655,29
1656,29
1657,29
1658,29
1659,29
1660,29
1661,29
1662,29
1663,29
1664,29
1665,29
1666,29
1667,29
1668,29
1669,29
1670,29
1671,29
1672,29
1673,29
1674,29
1675,29
1676,29
1677,29
1678,29
1679,29
1680,29
1681,29
1682,29
1683,29
1684,29
1685,29
1686,29
1687,29
1688,29
1689,29
1690,29
1691,29
1692,29
1693,29
1694,29
1695,29
1696,29
1697,29
1698,29
1699,29
1700,29
1701,29
1702,29
1703,29
1704,29
1705,29
1706,29
1707,29
1708,29
1709,29
1710,30
1711,30
1712,30
1713,30
1714,30
1715,30
1716,30
1717,30
1718,30
1719,30
1720,30
1721,30
1722,30
1723,30
1724,30
1725,30
1726,30
1727,30
1728,30
1729,30
1730,30
1731,30
1732,30
1733,30
1734,30
1735,30
1736,30
1737,30
1738,30
1739,30
1740,30
1741,30
1742,30
1743,30
1744,30
1745,30
1746,30
1747,30
1748,30
1749,30
1750,30
1751,30
1752,30
1753,30
1754,30
1755,30
1756,30
1757,30
1758,30
1759,30
1760,30
1761,30
1762,30
1763,30
1764,30
1765,30
1766,30
1767,31
1768,31
1769,31
1770,31
1771,31
1772,31
1773,31
1774,31
1775,31
1776,31
1777,31
1778,31
1779,31
1780,31
1781,31
1782,31
1783,31
1784,31
1785,31
1786,31
1787,31
1788,31
1789,31
1790,31
1791,31
1792,31
1793,31
1794,31
1795,31
1796,31
1797,31
1798,31
1799,31
1800,31
1801,31
1802,31
1803,31
1804,31
1805,31
1806,31
1807,31
1808,31
1809,31
1810,31
1811,31
1812,31
1813,31
1814,31
1815,31
1816,31
1817,31
1818,31
1819,31
1820,31
1821,31
1822,31
1823,31
1824,32
1825,32
1826,32
1827,32
1828,32
1829,32
1830,32
1831,32
1832,32
1833,32
1834,32
1835,32
1836,32
1837,32
1838,32
1839,32
1840,32
1841,32
1842,32
1843,32
1844,32
1845,32
1846,32
1847,32
1848,32
1849,32
1850,32
1851,32
1852,32
1853,32
1854,32
1855,32
1856,32
1857,32
1858,32
1859,32
1860,32
1861,32
1862,32
1863,32
1864,32
1865,32
1866,32
1867,32
1868,32
1869,32
1870,32
1871,32
1872,32
1873,32
1874,32
1875,32
1876,32
1877,32
1878,32
1879,32
1880,32
1881,33
1882,33
1883,33
1884,33
1885,33
1886,33
1887,33
1888,33
1889,33
1890,33
1891,33
1892,33
1893,33
1894,33
1895,33
1896,33
1897,33
1898,33
1899,33
1900,33
1901,33
1902,33
1903,33
1904,33
1905,33
1906,33
1907,33
1908,33
1909,33
1910,33
1911,33
1912,33
1913,33
1914,33
1915,33
1916,33
1917,33
1918,33
1919,33
1920,33
1921,33
1922,33
1923,33
1924,33
1925,33
1926,33
1927,33
1928,33
1929,33
1930,33
1931,33
1932,33
1933,33
1934,33
1935,33
1936,33
1937,33
1938,34
1939,34
1940,34
1941,34
1942,34
1943,34
1944,34
1945,34
1946,34
1947,34
1948,34
1949,34
1950,34
1951,34
1952,34
1953,34
1954,34
1955,34
1956,34
1957,34
1958,34
1959,34
1960,34
1961,34
1962,34
1963,34
1964,34
1965,34
1966,34
1967,34
1968,34
1969,34
1970,34
1971,34
1972,34
1973,34
1974,34
1975,34
1976,34
1977,34
1978,34
1979,34
1980,34
1981,34
1982,34
1983,34
1984,34
1985,34
1986,34
1987,34
1988,34
1989,34
1990,34
1991,34
1992,34
1993,34
1994,34
1995,35
1996,35
1997,35
1998,35
1999,35
2000,35
2001,35
2002,35
2003,35
2004,35
2005,35
2006,35
2007,35
2008,35
2009,35
2010,35
2011,35
2012,35
2013,35
2014,35
2015,35
2016,35
2017,35
2018,35
2019,35
2020,35
2021,35
2022,35
2023,35
2024,35
2025,35
2026,35
2027,35
2028,35
2029,35
2030,35
2031,35
2032,35
2033,35
2034,35
2035,35
2036,35
2037,35
2038,35
2039,35
2040,35
2041,35
2042,35
2043,35
2044,35
2045,35
2046,35
2047,35
2048,35
2049,35
2050,35
2051,35
2052,36
2053,36
2054,36
2055,36
2056,36
2057,36
2058,36
2059,36
2060,36
2061,36
2062,36
2063,36
2064,36
2065,36
2066,36
2067,36
2068,36
2069,36
2070,36
2071,36
2072,36
2073,36
2074,36
2075,36
2076,36
2077,36
2078,36
2079,36
2080,36
2081,36
2082,36
2083,36
2084,36
2085,36
2086,36
2087,36
2088,36
2089,36
2090,36
2091,36
2092,36
2093,36
2094,36
2095,36
2096,36
2097,36
2098,36
2099,36
2100,36
2101,36
2102,36
2103,36
2104,36
2105,36
2106,36
2107,36
2108,36
2109,37
2110,37
2111,37
2112,37
2113,37
2114,37
2115,37
2116,37
2117,37
2118,37
2119,37
2120,37
2121,37
2122,37
2123,37
2124,37
2125,37
2126,37
2127,37
2128,37
2129,37
2130,37
2131,37
2132,37
2133,37
2134,37
2135,37
2136,37
2137,37
2138,37
2139,37
2140,37
2141,37
2142,37
2143,37
2144,37
2145,37
2146,37
2147,37
2148,37
2149,37
2150,37
2151,37
2152,37
2153,37
2154,37
2155,37
2156,37
2157,37
2158,37
2159,37
2160,37
2161,37
2162,37
2163,37
2164,37
2165,37
2166,38
2167,38
2168,38
2169,38
2170,38
2171,38
2172,38
2173,38
2174,38
2175,38
2176,38
2177,38
2178,38
2179,38
2180,38
2181,38
2182,38
2183,38
2184,38
2185,38
2186,38
2187,38
2188,38
2189,38
2190,38
2191,38
2192,38
2193,38
2194,38
2195,38
2196,38
2197,38
2198,38
2199,38
2200,38
2201,38
2202,38
2203,38
2204,38
2205,38
2206,38
2207,38
2208,38
2209,38
2210,38
2211,38
2212,38
2213,38
2214,38
2215,38
2216,38
2217,38
2218,38
2219,38
2220,38
2221,38
2222,38
2223,39
2224,39
2225,39
2226,39
2227,39
2228,39
2229,39
2230,39
2231,39
2232,39
2233,39
2234,39
2235,39
2236,39
2237,39
2238,39
2239,39
2240,39
2241,39
2242,39
2243,39
2244,39
2245,39
2246,39
2247,39
2248,39
2249,39
2250,39
2251,39
2252,39
2253,39
2254,39
2255,39
2256,39
2257,39
2258,39
2259,39
2260,39
2261,39
2262,39
2263,39
2264,39
2265,39
2266,39
2267,39
2268,39
2269,39
2270,39
2271,39
2272,39
2273,39
2274,39
2275,39
2276,39
2277,39
2278,39
2279,39
2280,40
2281,40
2282,40
2283,40
2284,40
2285,40
2286,40
2287,40
2288,40
2289,40
2290,40
2291,40
2292,40
2293,40
2294,40
2295,40
2296,40
2297,40
2298,40
2299,40
2300,40
2301,40
2302,40
2303,40
2304,40
2305,40
2306,40
2307,40
2308,40
2309,40
2310,40
2311,40
2312,40
2313,40
2314,40
2315,40
2316,40
2317,40
2318,40
2319,40
2320,40
2321,40
2322,40
2323,40
2324,40
2325,40
2326,40
2327,40
2328,40
2329,40
2330,40
2331,40
2332,40
2333,40
2334,40
2335,40
2336,40
2337,41
2338,41
2339,41
2340,41
2341,41
2342,41
2343,41
2344,41
2345,41
2346,41
2347,41
2348,41
2349,41
2350,41
2351,41
2352,41
2353,41
2354,41
2355,41
2356,41
2357,41
2358,41
2359,41
2360,41
2361,41
2362,41
2363,41
2364,41
2365,41
2366,41
2367,41
2368,41
2369,41
2370,41
2371,41
2372,41
2373,41
2374,41
2375,41
2376,41
2377,41
2378,41
2379,41
2380,41
2381,41
2382,41
2383,41
2384,41
2385,41
2386,41
2387,41
2388,41
2389,41
2390,41
2391,41
2392,41
2393,41
2394,42
2395,42
2396,42
2397,42
2398,42
2399,42
2400,42
2401,42
2402,42
2403,42
2404,42
2405,42
2406,42
2407,42
2408,42
2409,42
2410,42
2411,42
2412,42
2413,42
2414,42
2415,42
2416,42
2417,42
2418,42
2419,42
2420,42
2421,42
2422,42
2423,42
2424,42
2425,42
2426,42
2427,42
2428,42
2429,42
2430,42
2431,42
2432,42
2433,42
2434,42
2435,42
2436,42
2437,42
2438,42
2439,42
2440,42
2441,42
2442,42
2443,42
2444,42
2445,42
2446,42
2447,42
2448,42
2449,42
2450,42
2451,43
2452,43
2453,43
2454,43
2455,43
2456,43
2457,43
2458,43
2459,43
2460,43
2461,43
2462,43
2463,43
2464,43
2465,43
2466,43
2467,43
2468,43
2469,43
2470,43
2471,43
2472,43
2473,43
2474,43
2475,43
2476,43
2477,43
2478,43
2479,43
2480,43
2481,43
2482,43
2483,43
2484,43
2485,43
2486,43
2487,43
2488,43
2489,43
2490,43
2491,43
2492,43
2493,43
2494,43
2495,43
2496,43
2497,43
2498,43
2499,43
2500,43
2501,43
2502,43
2503,43
2504,43
2505,43
2506,43
2507,43
2508,44
2509,44
2510,44
2511,44
2512,44
2513,44
2514,44
2515,44
2516,44
2517,44
2518,44
2519,44
2520,44
2521,44
2522,44
2523,44
2524,44
2525,44
2526,44
2527,44
2528,44
2529,44
2530,44
2531,44
2532,44
2533,44
2534,44
2535,44
2536,44
2537,44
2538,44
2539,44
2540,44
2541,44
2542,44
2543,44
2544,44
2545,44
2546,44
2547,44
2548,44
2549,44
2550,44
2551,44
2552,44
2553,44
2554,44
2555,44
2556,44
2557,44
2558,44
2559,44
2560,44
2561,44
2562,44
2563,44
2564,44
2565,45
2566,45
2567,45
2568,45
2569,45
2570,45
2571,45
2572,45
2573,45
2574,45
2575,45
2576,45
2577,45
2578,45
2579,45
2580,45
2581,45
2582,45
2583,45
2584,45
2585,45
2586,45
2587,45
2588,45
2589,45
2590,45
2591,45
2592,45
2593,45
2594,45
2595,45
2596,45
2597,45
2598,45
2599,45
2600,45
2601,45
2602,45
2603,45
2604,45
2605,45
2606,45
2607,45
2608,45
2609,45
2610,45
2611,45
2612,45
2613,45
2614,45
2615,45
2616,45
2617,45
2618,45
2619,45
2620,45
2621,45
2622,46
2623,46
2624,46
2625,46
2626,46
2627,46
2628,46
2629,46
2630,46
2631,46
2632,46
2633,46
2634,46
2635,46
2636,46
2637,46
2638,46
2639,46
2640,46
2641,46
2642,46
2643,46
2644,46
2645,46
2646,46
2647,46
2648,46
2649,46
2650,46
2651,46
2652,46
2653,46
2654,46
2655,46
2656,46
2657,46
2658,46
2659,46
2660,46
2661,46
2662,46
2663,46
2664,46
2665,46
2666,46
2667,46
2668,46
2669,46
2670,46
2671,46
2672,46
2673,46
2674,46
2675,46
2676,46
2677,46
2678,46
2679,47
2680,47
2681,47
2682,47
2683,47
2684,47
2685,47
2686,47
2687,47
2688,47
2689,47
2690,47
2691,47
2692,47
2693,47
2694,47
2695,47
2696,47
2697,47
2698,47
2699,47
2700,47
2701,47
2702,47
2703,47
2704,47
2705,47
2706,47
2707,47
2708,47
2709,47
2710,47
2711,47
2712,47
2713,47
2714,47
2715,47
2716,47
2717,47
2718,47
2719,47
2720,47
2721,47
2722,47
2723,47
2724,47
2725,47
2726,47
2727,47
2728,47
2729,47
2730,47
2731,47
2732,47
2733,47
2734,47
2735,47
2736,48
2737,48
2738,48
2739,48
2740,48
2741,48
2742,48
2743,48
2744,48
2745,48
2746,48
2747,48
2748,48
2749,48
2750,48
2751,48
2752,48
2753,48
2754,48
2755,48
2756,48
2757,48
2758,48
2759,48
2760,48
2761,48
2762,48
2763,48
2764,48
2765,48
2766,48
2767,48
2768,48
2769,48
2770,48
2771,48
2772,48
2773,48
2774,48
2775,48
2776,48
2777,48
2778,48
2779,48
2780,48
2781,48
2782,48
2783,48
2784,48
2785,48
2786,48
2787,48
2788,48
2789,48
2790,48
2791,48
2792,48
2793,48
2794,49
2795,49
2796,49
2797,49
2798,49
2799,49
2800,49
2801,49
2802,49
2803,49
2804,49
2805,49
2806,49
2807,49
2808,49
2809,49
2810,49
2811,49
2812,49
2813,49
2814,49
2815,49
2816,49
2817,49
2818,49
2819,49
2820,49
2821,49
2822,49
2823,49
2824,49
2825,49
2826,49
2827,49
2828,49
2829,49
2830,49
2831,49
2832,49
2833,49
2834,49
2835,49
2836,49
2837,49
2838,49
2839,49
2840,49
2841,49
2842,49
2843,49
2844,49
2845,49
2846,49
2847,49
2848,49
2849,49
2850,49
2851,49
2852,50
2853,50
2854,50
2855,50
2856,50
2857,50
2858,50
2859,50
2860,50
2861,50
2862,50
2863,50
2864,50
2865,50
2866,50
2867,50
2868,50
2869,50
2870,50
2871,50
2872,50
2873,50
2874,50
2875,50
2876,50
2877,50
2878,50
2879,50
2880,50
2881,50
2882,50
2883,50
2884,50
2885,50
2886,50
2887,50
2888,50
2889,50
2890,50
2891,50
2892,50
2893,50
2894,50
2895,50
2896,50
2897,50
2898,50
2899,50
2900,50
2901,50
2902,50
2903,50
2904,50
2905,50
2906,50
2907,50
2908,50
2909,50
2910,51
2911,51
2912,51
2913,51
2914,51
2915,51
2916,51
2917,51
2918,51
2919,51
2920,51
2921,51
2922,51
2923,51
2924,51
2925,51
2926,51
2927,51
2928,51
2929,51
2930,51
2931,51
2932,51
2933,51
2934,51
2935,51
2936,51
2937,51
2938,51
2939,51
2940,51
2941,51
2942,51
2943,51
2944,51
2945,51
2946,51
2947,51
2948,51
2949,51
2950,51
2951,51
2952,51
2953,51
2954,51
2955,51
2956,51
2957,51
2958,51
2959,51
2960,51
2961,51
2962,51
2963,51
2964,51
2965,51
2966,51
2967,51
2968,52
2969,52
2970,52
2971,52
2972,52
2973,52
2974,52
2975,52
2976,52
2977,52
2978,52
2979,52
2980,52
2981,52
2982,52
2983,52
2984,52
2985,52
2986,52
2987,52
2988,52
2989,52
2990,52
2991,52
2992,52
2993,52
2994,52
2995,52
2996,52
2997,52
2998,52
2999,52
3000,52
3001,52
3002,52
3003,52
3004,52
3005,52
3006,52
3007,52
3008,52
3009,52
3010,52
3011,52
3012,52
3013,52
3014,52
3015,52
3016,52
3017,52
3018,52
3019,52
3020,52
3021,52
3022,52
3023,52
3024,52
3025,52
3026,53
3027,53
3028,53
3029,53
3030,53
3031,53
3032,53
3033,53
3034,53
3035,53
3036,53
3037,53
3038,53
3039,53
3040,53
3041,53
3042,53
3043,53
3044,53
3045,53
3046,53
3047,53
3048,53
3049,53
3050,53
3051,53
3052,53
3053,53
3054,53
3055,53
3056,53
3057,53
3058,53
3059,53
3060,53
3061,53
3062,53
3063,53
3064,53
3065,53
3066,53
3067,53
3068,53
3069,53
3070,53
3071,53
3072,53
3073,53
3074,53
3075,53
3076,53
3077,53
3078,53
3079,53
3080,53
3081,53
3082,53
3083,53
3084,54
3085,54
3086,54
3087,54
3088,54
3089,54
3090,54
3091,54
3092,54
3093,54
3094,54
3095,54
3096,54
3097,54
3098,54
3099,54
3100,54
3101,54
3102,54
3103,54
3104,54
3105,54
3106,54
3107,54
3108,54
3109,54
3110,54
3111,54
3112,54
3113,54
3114,54
3115,54
3116,54
3117,54
3118,54
3119,54
3120,54
3121,54
3122,54
3123,54
3124,54
3125,54
3126,54
3127,54
3128,54
3129,54
3130,54
3131,54
3132,54
3133,54
3134,54
3135,54
3136,54
3137,54
3138,54
3139,54
3140,54
3141,54
3142,55
3143,55
3144,55
3145,55
3146,55
3147,55
3148,55
3149,55
3150,55
3151,55
3152,55
3153,55
3154,55
3155,55
3156,55
3157,55
3158,55
3159,55
3160,55
3161,55
3162,55
3163,55
3164,55
3165,55
3166,55
3167,55
3168,55
3169,55
3170,55
3171,55
3172,55
3173,55
3174,55
3175,55
3176,55
3177,55
3178,55
3179,55
3180,55
3181,55
3182,55
3183,55
3184,55
3185,55
3186,55
3187,55
3188,55
3189,55
3190,55
3191,55
3192,55
3193,55
3194,55
3195,55
3196,55
3197,55
3198,55
3199,55
3200,56
3201,56
3202,56
3203,56
3204,56
3205,56
3206,56
3207,56
3208,56
3209,56
3210,56
3211,56
3212,56
3213,56
3214,56
3215,56
3216,56
3217,56
3218,56
3219,56
3220,56
3221,56
3222,56
3223,56
3224,56
3225,56
3226,56
3227,56
3228,56
3229,56
3230,56
3231,56
3232,56
3233,56
3234,56
3235,56
3236,56
3237,56
3238,56
3239,56
3240,56
3241,56
3242,56
3243,56
3244,56
3245,56
3246,56
3247,56
3248,56
3249,56
3250,56
3251,56
3252,56
3253,56
3254,56
3255,56
3256,56
3257,56
3258,57
3259,57
3260,57
3261,57
3262,57
3263,57
3264,57
3265,57
3266,57
3267,57
3268,57
3269,57
3270,57
3271,57
3272,57
3273,57
3274,57
3275,57
3276,57
3277,57
3278,57
3279,57
3280,57
3281,57
3282,57
3283,57
3284,57
3285,57
3286,57
3287,57
3288,57
3289,57
3290,57
3291,57
3292,57
3293,57
3294,57
3295,57
3296,57
3297,57
3298,57
3299,57
3300,57
3301,57
3302,57
3303,57
3304,57
3305,57
3306,57
3307,57
3308,57
3309,57
3310,57
3311,57
3312,57
3313,57
3314,57
3315,57
3316,58
3317,58
3318,58
3319,58
3320,58
3321,58
3322,58
3323,58
3324,58
3325,58
3326,58
3327,58
3328,58
3329,58
3330,58
3331,58
3332,58
3333,58
3334,58
3335,58
3336,58
3337,58
3338,58
3339,58
3340,58
3341,58
3342,58
3343,58
3344,58
3345,58
3346,58
3347,58
3348,58
3349,58
3350,58
3351,58
3352,58
3353,58
3354,58
3355,58
3356,58
3357,58
3358,58
3359,58
3360,58
3361,58
3362,58
3363,58
3364,58
3365,58
3366,58
3367,58
3368,58
3369,58
3370,58
3371,58
3372,58
3373,58
3374,59
3375,59
3376,59
3377,59
3378,59
3379,59
3380,59
3381,59
3382,59
3383,59
3384,59
3385,59
3386,59
3387,59
3388,59
3389,59
3390,59
3391,59
3392,59
3393,59
3394,59
3395,59
3396,59
3397,59
3398,59
3399,59
3400,59
3401,59
3402,59
3403,59
3404,59
3405,59
3406,59
3407,59
3408,59
3409,59
3410,59
3411,59
3412,59
3413,59
3414,59
3415,59
3416,59
3417,59
3418,59
3419,59
3420,59
3421,59
3422,59
3423,59
3424,59
3425,59
3426,59
3427,59
3428,59
3429,59
3430,59
3431,59
3432,60
3433,60
3434,60
3435,60
3436,60
3437,60
3438,60
3439,60
3440,60
3441,60
3442,60
3443,60
3444,60
3445,60
3446,60
3447,60
3448,60
3449,60
3450,60
3451,60
3452,60
3453,60
3454,60
3455,60
3456,60
3457,60
3458,60
3459,60
3460,60
3461,60
3462,60
3463,60
3464,60
3465,60
3466,60
3467,60
3468,60
3469,60
3470,60
3471,60
3472,60
3473,60
3474,60
3475,60
3476,60
3477,60
3478,60
3479,60
3480,60
3481,60
3482,60
3483,60
3484,60
3485,60
3486,60
3487,60
3488,60
3489,60
3490,61
3491,61
3492,61
3493,61
3494,61
3495,61
3496,61
3497,61
3498,61
3499,61
3500,61
3501,61
3502,61
3503,61
3504,61
3505,61
3506,61
3507,61
3508,61
3509,61
3510,61
3511,61
3512,61
3513,61
3514,61
3515,61
3516,61
3517,61
3518,61
3519,61
3520,61
3521,61
3522,61
3523,61
3524,61
3525,61
3526,61
3527,61
3528,61
3529,61
3530,61
3531,61
3532,61
3533,61
3534,61
3535,61
3536,61
3537,61
3538,61
3539,61
3540,61
3541,61
3542,61
3543,61
3544,61
3545,61
3546,61
3547,61
3548,62
3549,62
3550,62
3551,62
3552,62
3553,62
3554,62
3555,62
3556,62
3557,62
3558,62
3559,62
3560,62
3561,62
3562,62
3563,62
3564,62
3565,62
3566,62
3567,62
3568,62
3569,62
3570,62
3571,62
3572,62
3573,62
3574,62
3575,62
3576,62
3577,62
3578,62
3579,62
3580,62
3581,62
3582,62
3583,62
3584,62
3585,62
3586,62
3587,62
3588,62
3589,62
3590,62
3591,62
3592,62
3593,62
3594,62
3595,62
3596,62
3597,62
3598,62
3599,62
3600,62
3601,62
3602,62
3603,62
3604,62
3605,62
3606,63
3607,63
3608,63
3609,63
3610,63
3611,63
3612,63
3613,63
3614,63
3615,63
3616,63
3617,63
3618,63
3619,63
3620,63
3621,63
3622,63
3623,63
3624,63
3625,63
3626,63
3627,63
3628,63
3629,63
3630,63
3631,63
3632,63
3633,63
3634,63
3635,63
3636,63
3637,63
3638,63
3639,63
3640,63
3641,63
3642,63
3643,63
3644,63
3645,63
3646,63
3647,63
3648,63
3649,63
3650,63
3651,63
3652,63
3653,63
3654,63
3655,63
3656,63
3657,63
3658,63
3659,63
3660,63
3661,63
3662,63
3663,63
3664,64
3665,64
3666,64
3667,64
3668,64
3669,64
3670,64
3671,64
3672,64
3673,64
3674,64
3675,64
3676,64
3677,64
3678,64
3679,64
3680,64
3681,64
3682,64
3683,64
3684,64
3685,64
3686,64
3687,64
3688,64
3689,64
3690,64
3691,64
3692,64
3693,64
3694,64
3695,64
3696,64
3697,64
3698,64
3699,64
3700,64
3701,64
3702,64
3703,64
3704,64
3705,64
3706,64
3707,64
3708,64
3709,64
3710,64
3711,64
3712,64
3713,64
3714,64
3715,64
3716,64
3717,64
3718,64
3719,64
3720,64
3721,64
3722,65
3723,65
3724,65
3725,65
3726,65
3727,65
3728,65
3729,65
3730,65
3731,65
3732,65
3733,65
3734,65
3735,65
3736,65
3737,65
3738,65
3739,65
3740,65
3741,65
3742,65
3743,65
3744,65
3745,65
3746,65
3747,65
3748,65
3749,65
3750,65
3751,65
3752,65
3753,65
3754,65
3755,65
3756,65
3757,65
3758,65
3759,65
3760,65
3761,65
3762,65
3763,65
3764,65
3765,65
3766,65
3767,65
3768,65
3769,65
3770,65
3771,65
3772,65
3773,65
3774,65
3775,65
3776,65
3777,65
3778,65
3779,65
3780,66
3781,66
3782,66
3783,66
3784,66
3785,66
3786,66
3787,66
3788,66
3789,66
3790,66
3791,66
3792,66
3793,66
3794,66
3795,66
3796,66
3797,66
3798,66
3799,66
3800,66
3801,66
3802,66
3803,66
3804,66
3805,66
3806,66
3807,66
3808,66
3809,66
3810,66
3811,66
3812,66
3813,66
3814,66
3815,66
3816,66
3817,66
3818,66
3819,66
3820,66
3821,66
3822,66
3823,66
3824,66
3825,66
3826,66
3827,66
3828,66
3829,66
3830,66
3831,66
3832,66
3833,66
3834,66
3835,66
3836,66
3837,66
3838,67
3839,67
3840,67
3841,67
3842,67
3843,67
3844,67
3845,67
3846,67
3847,67
3848,67
3849,67
3850,67
3851,67
3852,67
3853,67
3854,67
3855,67
3856,67
3857,67
3858,67
3859,67
3860,67
3861,67
3862,67
3863,67
3864,67
3865,67
3866,67
3867,67
3868,67
3869,67
3870,67
3871,67
3872,67
3873,67
3874,67
3875,67
3876,67
3877,67
3878,67
3879,67
3880,67
3881,67
3882,67
3883,67
3884,67
3885,67
3886,67
3887,67
3888,67
3889,67
3890,67
3891,67
3892,67
3893,67
3894,67
3895,67
3896,68
3897,68
3898,68
3899,68
3900,68
3901,68
3902,68
3903,68
3904,68
3905,68
3906,68
3907,68
3908,68
3909,68
3910,68
3911,68
3912,68
3913,68
3914,68
3915,68
3916,68
3917,68
3918,68
3919,68
3920,68
3921,68
3922,68
3923,68
3924,68
3925,68
3926,68
3927,68
3928,68
3929,68
3930,68
3931,68
3932,68
3933,68
3934,68
3935,68
3936,68
3937,68
3938,68
3939,68
3940,68
3941,68
3942,68
3943,68
3944,68
3945,68
3946,68
3947,68
3948,68
3949,68
3950,68
3951,68
3952,68
3953,68
3954,69
3955,69
3956,69
3957,69
3958,69
3959,69
3960,69
3961,69
3962,69
3963,69
3964,69
3965,69
3966,69
3967,69
3968,69
3969,69
3970,69
3971,69
3972,69
3973,69
3974,69
3975,69
3976,69
3977,69
3978,69
3979,69
3980,69
3981,69
3982,69
3983,69
3984,69
3985,69
3986,69
3987,69
3988,69
3989,69
3990,69
3991,69
3992,69
3993,69
3994,69
3995,69
3996,69
3997,69
3998,69
3999,69
4000,69
4001,69
4002,69
4003,69
4004,69
4005,69
4006,69
4007,69
4008,69
4009,69
4010,69
4011,69
4012,70
4013,70
4014,70
4015,70
4016,70
4017,70
4018,70
4019,70
4020,70
4021,70
4022,70
4023,70
4024,70
4025,70
4026,70
4027,70
4028,70
4029,70
4030,70
4031,70
4032,70
4033,70
4034,70
4035,70
4036,70
4037,70
4038,70
4039,70
4040,70
4041,70
4042,70
4043,70
4044,70
4045,70
4046,70
4047,70
4048,70
4049,70
4050,70
4051,70
4052,70
4053,70
4054,70
4055,70
4056,70
4057,70
4058,70
4059,70
4060,70
4061,70
4062,70
4063,70
4064,70
4065,70
4066,70
4067,70
4068,70
4069,70
4070,71
4071,71
4072,71
4073,71
4074,71
4075,71
4076,71
4077,71
4078,71
4079,71
4080,71
4081,71
4082,71
4083,71
4084,71
4085,71
4086,71
4087,71
4088,71
4089,71
4090,71
4091,71
4092,71
4093,71
4094,71
4095,71
4096,71
4097,71
4098,71
4099,71
4100,71
4101,71
4102,71
4103,71
4104,71
4105,71
4106,71
4107,71
4108,71
4109,71
4110,71
4111,71
4112,71
4113,71
4114,71
4115,71
4116,71
4117,71
4118,71
4119,71
4120,71
4121,71
4122,71
4123,71
4124,71
4125,71
4126,71
4127,71
4128,72
4129,72
4130,72
4131,72
4132,72
4133,72
4134,72
4135,72
4136,72
4137,72
4138,72
4139,72
4140,72
4141,72
4142,72
4143,72
4144,72
4145,72
4146,72
4147,72
4148,72
4149,72
4150,72
4151,72
4152,72
4153,72
4154,72
4155,72
4156,72
4157,72
4158,72
4159,72
4160,72
4161,72
4162,72
4163,72
4164,72
4165,72
4166,72
4167,72
4168,72
4169,72
4170,72
4171,72
4172,72
4173,72
4174,72
4175,72
4176,72
4177,72
4178,72
4179,72
4180,72
4181,72
4182,72
4183,72
4184,72
4185,72
4186,73
4187,73
4188,73
4189,73
4190,73
4191,73
4192,73
4193,73
4194,73
4195,73
4196,73
4197,73
4198,73
4199,73
4200,73
4201,73
4202,73
4203,73
4204,73
4205,73
4206,73
4207,73
4208,73
4209,73
4210,73
4211,73
4212,73
4213,73
4214,73
4215,73
4216,73
4217,73
4218,73
4219,73
4220,73
4221,73
4222,73
4223,73
4224,73
4225,73
4226,73
4227,73
4228,73
4229,73
4230,73
4231,73
4232,73
4233,73
4234,73
4235,73
4236,73
4237,73
4238,73
4239,73
4240,73
4241,73
4242,73
4243,73
4244,74
4245,74
4246,74
4247,74
4248,74
4249,74
4250,74
4251,74
4252,74
4253,74
4254,74
4255,74
4256,74
4257,74
4258,74
4259,74
4260,74
4261,74
4262,74
4263,74
4264,74
4265,74
4266,74
4267,74
4268,74
4269,74
4270,74
4271,74
4272,74
4273,74
4274,74
4275,74
4276,74
4277,74
4278,74
4279,74
4280,74
4281,74
4282,74
4283,74
4284,74
4285,74
4286,74
4287,74
4288,74
4289,74
4290,74
4291,74
4292,74
4293,74
4294,74
4295,74
4296,74
4297,74
4298,74
4299,74
4300,74
4301,74
4302,75
4303,75
4304,75
4305,75
4306,75
4307,75
4308,75
4309,75
4310,75
4311,75
4312,75
4313,75
4314,75
4315,75
4316,75
4317,75
4318,75
4319,75
4320,75
4321,75
4322,75
4323,75
4324,75
4325,75
4326,75
4327,75
4328,75
4329,75
4330,75
4331,75
4332,75
4333,75
4334,75
4335,75
4336,75
4337,75
4338,75
4339,75
4340,75
4341,75
4342,75
4343,75
4344,75
4345,75
4346,75
4347,75
4348,75
4349,75
4350,75
4351,75
4352,75
4353,75
4354,75
4355,75
4356,75
4357,75
4358,75
4359,75
4360,76
4361,76
4362,76
4363,76
4364,76
4365,76
4366,76
4367,76
4368,76
4369,76
4370,76
4371,76
4372,76
4373,76
4374,76
4375,76
4376,76
4377,76
4378,76
4379,76
4380,76
4381,76
4382,76
4383,76
4384,76
4385,76
4386,76
4387,76
4388,76
4389,76
4390,76
4391,76
4392,76
4393,76
4394,76
4395,76
4396,76
4397,76
4398,76
4399,76
4400,76
4401,76
4402,76
4403,76
4404,76
4405,76
4406,76
4407,76
4408,76
4409,76
4410,76
4411,76
4412,76
4413,76
4414,76
4415,76
4416,76
4417,76
4418,77
4419,77
4420,77
4421,77
4422,77
4423,77
4424,77
4425,77
4426,77
4427,77
4428,77
4429,77
4430,77
4431,77
4432,77
4433,77
4434,77
4435,77
4436,77
4437,77
4438,77
4439,77
4440,77
4441,77
4442,77
4443,77
4444,77
4445,77
4446,77
4447,77
4448,77
4449,77
4450,77
4451,77
4452,77
4453,77
4454,77
4455,77
4456,77
4457,77
4458,77
4459,77
4460,77
4461,77
4462,77
4463,77
4464,77
4465,77
4466,77
4467,77
4468,77
4469,77
4470,77
4471,77
4472,77
4473,77
4474,77
4475,77
4476,78
4477,78
4478,78
4479,78
4480,78
4481,78
4482,78
4483,78
4484,78
4485,78
4486,78
4487,78
4488,78
4489,78
4490,78
4491,78
4492,78
4493,78
4494,78
4495,78
4496,78
4497,78
4498,78
4499,78
4500,78
4501,78
4502,78
4503,78
4504,78
4505,78
4506,78
4507,78
4508,78
4509,78
4510,78
4511,78
4512,78
4513,78
4514,78
4515,78
4516,78
4517,78
4518,78
4519,78
4520,78
4521,78
4522,78
4523,78
4524,78
4525,78
4526,78
4527,78
4528,78
4529,78
4530,78
4531,78
4532,78
4533,78
4534,79
4535,79
4536,79
4537,79
4538,79
4539,79
4540,79
4541,79
4542,79
4543,79
4544,79
4545,79
4546,79
4547,79
4548,79
4549,79
4550,79
4551,79
4552,79
4553,79
4554,79
4555,79
4556,79
4557,79
4558,79
4559,79
4560,79
4561,79
4562,79
4563,79
4564,79
4565,79
4566,79
4567,79
4568,79
4569,79
4570,79
4571,79
4572,79
4573,79
4574,79
4575,79
4576,79
4577,79
4578,79
4579,79
4580,79
4581,79
4582,79
4583,79
4584,79
4585,79
4586,79
4587,79
4588,79
4589,79
4590,79
4591,79
4592,80
4593,80
4594,80
4595,80
4596,80
4597,80
4598,80
4599,80
4600,80
4601,80
4602,80
4603,80
4604,80
4605,80
4606,80
4607,80
4608,80
4609,80
4610,80
4611,80
4612,80
4613,80
4614,80
4615,80
4616,80
4617,80
4618,80
4619,80
4620,80
4621,80
4622,80
4623,80
4624,80
4625,80
4626,80
4627,80
4628,80
4629,80
4630,80
4631,80
4632,80
4633,80
4634,80
4635,80
4636,80
4637,80
4638,80
4639,80
4640,80
4641,80
4642,80
4643,80
4644,80
4645,80
4646,80
4647,80
4648,80
4649,80
4650,81
4651,81
4652,81
4653,81
4654,81
4655,81
4656,81
4657,81
4658,81
4659,81
4660,81
4661,81
4662,81
4663,81
4664,81
4665,81
4666,81
4667,81
4668,81
4669,81
4670,81
4671,81
4672,81
4673,81
4674,81
4675,81
4676,81
4677,81
4678,81
4679,81
4680,81
4681,81
4682,81
4683,81
4684,81
4685,81
4686,81
4687,81
4688,81
4689,81
4690,81
4691,81
4692,81
4693,81
4694,81
4695,81
4696,81
4697,81
4698,81
4699,81
4700,81
4701,81
4702,81
4703,81
4704,81
4705,81
4706,81
4707,81
4708,82
4709,82
4710,82
4711,82
4712,82
4713,82
4714,82
4715,82
4716,82
4717,82
4718,82
4719,82
4720,82
4721,82
4722,82
4723,82
4724,82
4725,82
4726,82
4727,82
4728,82
4729,82
4730,82
4731,82
4732,82
4733,82
4734,82
4735,82
4736,82
4737,82
4738,82
4739,82
4740,82
4741,82
4742,82
4743,82
4744,82
4745,82
4746,82
4747,82
4748,82
4749,82
4750,82
4751,82
4752,82
4753,82
4754,82
4755,82
4756,82
4757,82
4758,82
4759,82
4760,82
4761,82
4762,82
4763,82
4764,82
4765,82
4766,83
4767,83
4768,83
4769,83
4770,83
4771,83
4772,83
4773,83
4774,83
4775,83
4776,83
4777,83
4778,83
4779,83
4780,83
4781,83
4782,83
4783,83
4784,83
4785,83
4786,83
4787,83
4788,83
4789,83
4790,83
4791,83
4792,83
4793,83
4794,83
4795,83
4796,83
4797,83
4798,83
4799,83
4800,83
4801,83
4802,83
4803,83
4804,83
4805,83
4806,83
4807,83
4808,83
4809,83
4810,83
4811,83
4812,83
4813,83
4814,83
4815,83
4816,83
4817,83
4818,83
4819,83
4820,83
4821,83
4822,83
4823,83
4824,84
4825,84
4826,84
4827,84
4828,84
4829,84
4830,84
4831,84
4832,84
4833,84
4834,84
4835,84
4836,84
4837,84
4838,84
4839,84
4840,84
4841,84
4842,84
4843,84
4844,84
4845,84
4846,84
4847,84
4848,84
4849,84
4850,84
4851,84
4852,84
4853,84
4854,84
4855,84
4856,84
4857,84
4858,84
4859,84
4860,84
4861,84
4862,84
4863,84
4864,84
4865,84
4866,84
4867,84
4868,84
4869,84
4870,84
4871,84
4872,84
4873,84
4874,84
4875,84
4876,84
4877,84
4878,84
4879,84
4880,84
4881,84
4882,85
4883,85
4884,85
4885,85
4886,85
4887,85
4888,85
4889,85
4890,85
4891,85
4892,85
4893,85
4894,85
4895,85
4896,85
4897,85
4898,85
4899,85
4900,85
4901,85
4902,85
4903,85
4904,85
4905,85
4906,85
4907,85
4908,85
4909,85
4910,85
4911,85
4912,85
4913,85
4914,85
4915,85
4916,85
4917,85
4918,85
4919,85
4920,85
4921,85
4922,85
4923,85
4924,85
4925,85
4926,85
4927,85
4928,85
4929,85
4930,85
4931,85
4932,85
4933,85
4934,85
4935,85
4936,85
4937,85
4938,85
4939,85
4940,86
4941,86
4942,86
4943,86
4944,86
4945,86
4946,86
4947,86
4948,86
4949,86
4950,86
4951,86
4952,86
4953,86
4954,86
4955,86
4956,86
4957,86
4958,86
4959,86
4960,86
4961,86
4962,86
4963,86
4964,86
4965,86
4966,86
4967,86
4968,86
4969,86
4970,86
4971,86
4972,86
4973,86
4974,86
4975,86
4976,86
4977,86
4978,86
4979,86
4980,86
4981,86
4982,86
4983,86
4984,86
4985,86
4986,86
4987,86
4988,86
4989,86
4990,86
4991,86
4992,86
4993,86
4994,86
4995,86
4996,86
4997,86
4998,87
4999,87
5000,87
5001,87
5002,87
5003,87
5004,87
5005,87
5006,87
5007,87
5008,87
5009,87
5010,87
5011,87
5012,87
5013,87
5014,87
5015,87
5016,87
5017,87
5018,87
5019,87
5020,87
5021,87
5022,87
5023,87
5024,87
5025,87
5026,87
5027,87
5028,87
5029,87
5030,87
5031,87
5032,87
5033,87
5034,87
5035,87
5036,87
5037,87
5038,87
5039,87
5040,87
5041,87
5042,87
5043,87
5044,87
5045,87
5046,87
5047,87
5048,87
5049,87
5050,87
5051,87
5052,87
5053,87
5054,87
5055,87
5056,88
5057,88
5058,88
5059,88
5060,88
5061,88
5062,88
5063,88
5064,88
5065,88
5066,88
5067,88
5068,88
5069,88
5070,88
5071,88
5072,88
5073,88
5074,88
5075,88
5076,88
5077,88
5078,88
5079,88
5080,88
5081,88
5082,88
5083,88
5084,88
5085,88
5086,88
5087,88
5088,88
5089,88
5090,88
5091,88
5092,88
5093,88
5094,88
5095,88
5096,88
5097,88
5098,88
5099,88
5100,88
5101,88
5102,88
5103,88
5104,88
5105,88
5106,88
5107,88
5108,88
5109,88
5110,88
5111,88
5112,88
5113,88
5114,89
5115,89
5116,89
5117,89
5118,89
5119,89
5120,89
5121,89
5122,89
5123,89
5124,89
5125,89
5126,89
5127,89
5128,89
5129,89
5130,89
5131,89
5132,89
5133,89
5134,89
5135,89
5136,89
5137,89
5138,89
5139,89
5140,89
5141,89
5142,89
5143,89
5144,89
5145,89
5146,89
5147,89
5148,89
5149,89
5150,89
5151,89
5152,89
5153,89
5154,89
5155,89
5156,89
5157,89
5158,89
5159,89
5160,89
5161,89
5162,89
5163,89
5164,89
5165,89
5166,89
5167,89
5168,89
5169,89
5170,89
5171,89
5172,90
5173,90
5174,90
5175,90
5176,90
5177,90
5178,90
5179,90
5180,90
5181,90
5182,90
5183,90
5184,90
5185,90
5186,90
5187,90
5188,90
5189,90
5190,90
5191,90
5192,90
5193,90
5194,90
5195,90
5196,90
5197,90
5198,90
5199,90
5200,90
5201,90
5202,90
5203,90
5204,90
5205,90
5206,90
5207,90
5208,90
5209,90
5210,90
5211,90
5212,90
5213,90
5214,90
5215,90
5216,90
5217,90
5218,90
5219,90
5220,90
5221,90
5222,90
5223,90
5224,90
5225,90
5226,90
5227,90
5228,90
5229,90
5230,91
5231,91
5232,91
5233,91
5234,91
5235,91
5236,91
5237,91
5238,91
5239,91
5240,91
5241,91
5242,91
5243,91
5244,91
5245,91
5246,91
5247,91
5248,91
5249,91
5250,91
5251,91
5252,91
5253,91
5254,91
5255,91
5256,91
5257,91
5258,91
5259,91
5260,91
5261,91
5262,91
5263,91
5264,91
5265,91
5266,91
5267,91
5268,91
5269,91
5270,91
5271,91
5272,91
5273,91
5274,91
5275,91
5276,91
5277,91
5278,91
5279,91
5280,91
5281,91
5282,91
5283,91
5284,91
5285,91
5286,91
5287,91
5288,92
5289,92
5290,92
5291,92
5292,92
5293,92
5294,92
5295,92
5296,92
5297,92
5298,92
5299,92
5300,92
5301,92
5302,92
5303,92
5304,92
5305,92
5306,92
5307,92
5308,92
5309,92
5310,92
5311,92
5312,92
5313,92
5314,92
5315,92
5316,92
5317,92
5318,92
5319,92
5320,92
5321,92
5322,92
5323,92
5324,92
5325,92
5326,92
5327,92
5328,92
5329,92
5330,92
5331,92
5332,92
5333,92
5334,92
5335,92
5336,92
5337,92
5338,92
5339,92
5340,92
5341,92
5342,92
5343,92
5344,92
5345,92
5346,93
5347,93
5348,93
5349,93
5350,93
5351,93
5352,93
5353,93
5354,93
5355,93
5356,93
5357,93
5358,93
5359,93
5360,93
5361,93
5362,93
5363,93
5364,93
5365,93
5366,93
5367,93
5368,93
5369,93
5370,93
5371,93
5372,93
5373,93
5374,93
5375,93
5376,93
5377,93
5378,93
5379,93
5380,93
5381,93
5382,93
5383,93
5384,93
5385,93
5386,93
5387,93
5388,93
5389,93
5390,93
5391,93
5392,93
5393,93
5394,93
5395,93
5396,93
5397,93
5398,93
5399,93
5400,93
5401,93
5402,93
5403,93
5404,94
5405,94
5406,94
5407,94
5408,94
5409,94
5410,94
5411,94
5412,94
5413,94
5414,94
5415,94
5416,94
5417,94
5418,94
5419,94
5420,94
5421,94
5422,94
5423,94
5424,94
5425,94
5426,94
5427,94
5428,94
5429,94
5430,94
5431,94
5432,94
5433,94
5434,94
5435,94
5436,94
5437,94
5438,94
5439,94
5440,94
5441,94
5442,94
5443,94
5444,94
5445,94
5446,94
5447,94
5448,94
5449,94
5450,94
5451,94
5452,94
5453,94
5454,94
5455,94
5456,94
5457,94
5458,94
5459,94
5460,94
5461,94
5462,95
5463,95
5464,95
5465,95
5466,95
5467,95
5468,95
5469,95
5470,95
5471,95
5472,95
5473,95
5474,95
5475,95
5476,95
5477,95
5478,95
5479,95
5480,95
5481,95
5482,95
5483,95
5484,95
5485,95
5486,95
5487,95
5488,95
5489,95
5490,95
5491,95
5492,95
5493,95
5494,95
5495,95
5496,95
5497,95
5498,95
5499,95
5500,95
5501,95
5502,95
5503,95
5504,95
5505,95
5506,95
5507,95
5508,95
5509,95
5510,95
5511,95
5512,95
5513,95
5514,95
5515,95
5516,95
5517,95
5518,95
5519,95
5520,96
5521,96
5522,96
5523,96
5524,96
5525,96
5526,96
5527,96
5528,96
5529,96
5530,96
5531,96
5532,96
5533,96
5534,96
5535,96
5536,96
5537,96
5538,96
5539,96
5540,96
5541,96
5542,96
5543,96
5544,96
5545,96
5546,96
5547,96
5548,96
5549,96
5550,96
5551,96
5552,96
5553,96
5554,96
5555,96
5556,96
5557,96
5558,96
5559,96
5560,96
5561,96
5562,96
5563,96
5564,96
5565,96
5566,96
5567,96
5568,96
5569,96
5570,96
5571,96
5572,96
5573,96
5574,96
5575,96
5576,96
5577,96
5578,97
5579,97
5580,97
5581,97
5582,97
5583,97
5584,97
5585,97
5586,97
5587,97
5588,97
5589,97
5590,97
5591,97
5592,97
5593,97
5594,97
5595,97
5596,97
5597,97
5598,97
5599,97
5600,97
5601,97
5602,97
5603,97
5604,97
5605,97
5606,97
5607,97
5608,97
5609,97
5610,97
5611,97
5612,97
5613,97
5614,97
5615,97
5616,97
5617,97
5618,97
5619,97
5620,97
5621,97
5622,97
5623,97
5624,97
5625,97
5626,97
5627,97
5628,97
5629,97
5630,97
5631,97
5632,97
5633,97
5634,97
5635,97
5636,98
5637,98
5638,98
5639,98
5640,98
5641,98
5642,98
5643,98
5644,98
5645,98
5646,98
5647,98
5648,98
5649,98
5650,98
5651,98
5652,98
5653,98
5654,98
5655,98
5656,98
5657,98
5658,98
5659,98
5660,98
5661,98
5662,98
5663,98
5664,98
5665,98
5666,98
5667,98
5668,98
5669,98
5670,98
5671,98
5672,98
5673,98
5674,98
5675,98
5676,98
5677,98
5678,98
5679,98
5680,98
5681,98
5682,98
5683,98
5684,98
5685,98
5686,98
5687,98
5688,98
5689,98
5690,98
5691,98
5692,98
5693,98
5694,99
5695,99
5696,99
5697,99
5698,99
5699,99
5700,99
5701,99
5702,99
5703,99
5704,99
5705,99
5706,99
5707,99
5708,99
5709,99
5710,99
5711,99
5712,99
5713,99
5714,99
5715,99
5716,99
5717,99
5718,99
5719,99
5720,99
5721,99
5722,99
5723,99
5724,99
5725,99
5726,99
5727,99
5728,99
5729,99
5730,99
5731,99
5732,99
5733,99
5734,99
5735,99
5736,99
5737,99
5738,99
5739,99
5740,99
5741,99
5742,99
5743,99
5744,99
5745,99
5746,99
5747,99
5748,99
5749,99
5750,99
5751,99
5752,100
5753,100
5754,100
5755,100
5756,100
5757,100
5758,100
5759,100
5760,100
5761,100
5762,100
5763,100
5764,100
5765,100
5766,100
5767,100
5768,100
5769,100
5770,100
5771,100
5772,100
5773,100
5774,100
5775,100
5776,100
5777,100
5778,100
5779,100
5780,100
5781,100
5782,100
5783,100
5784,100
5785,100
5786,100
5787,100
5788,100
5789,100
5790,100
5791,100
5792,100
5793,100
5794,100
5795,100
5796,100
5797,100
5798,100
5799,100
5800,100
5801,100
5802,100
5803,100
5804,100
5805,100
5806,100
5807,100
5808,100
5809,100
5810,101
5811,101
5812,101
5813,101
5814,101
5815,101
5816,101
5817,101
5818,101
5819,101
5820,101
5821,101
5822,101
5823,101
5824,101
5825,101
5826,101
5827,101
5828,101
5829,101
5830,101
5831,101
5832,101
5833,101
5834,101
5835,101
5836,101
5837,101
5838,101
5839,101
5840,101
5841,101
5842,101
5843,101
5844,101
5845,101
5846,101
5847,101
5848,101
5849,101
5850,101
5851,101
5852,101
5853,101
5854,101
5855,101
5856,101
5857,101
5858,101
5859,101
5860,101
5861,101
5862,101
5863,101
5864,101
5865,101
5866,101
5867,101
5868,102
5869,102
5870,102
5871,102
5872,102
5873,102
5874,102
5875,102
5876,102
5877,102
5878,102
5879,102
5880,102
5881,102
5882,102
5883,102
5884,102
5885,102
5886,102
5887,102
5888,102
5889,102
5890,102
5891,102
5892,102
5893,102
5894,102
5895,102
5896,102
5897,102
5898,102
5899,102
5900,102
5901,102
5902,102
5903,102
5904,102
5905,102
5906,102
5907,102
5908,102
5909,102
5910,102
5911,102
5912,102
5913,102
5914,102
5915,102
5916,102
5917,102
5918,102
5919,102
5920,102
5921,102
5922,102
5923,102
5924,102
5925,102
5926,103
5927,103
5928,103
5929,103
5930,103
5931,103
5932,103
5933,103
5934,103
5935,103
5936,103
5937,103
5938,103
5939,103
5940,103
5941,103
5942,103
5943,103
5944,103
5945,103
5946,103
5947,103
5948,103
5949,103
5950,103
5951,103
5952,103
5953,103
5954,103
5955,103
5956,103
5957,103
5958,103
5959,103
5960,103
5961,103
5962,103
5963,103
5964,103
5965,103
5966,103
5967,103
5968,103
5969,103
5970,103
5971,103
5972,103
5973,103
5974,103
5975,103
5976,103
5977,103
5978,103
5979,103
5980,103
5981,103
5982,103
5983,103
5984,104
5985,104
5986,104
5987,104
5988,104
5989,104
5990,104
5991,104
5992,104
5993,104
5994,104
5995,104
5996,104
5997,104
5998,104
5999,104
6000,104
6001,104
6002,104
6003,104
6004,104
6005,104
6006,104
6007,104
6008,104
6009,104
6010,104
6011,104
6012,104
6013,104
6014,104
6015,104
6016,104
6017,104
6018,104
6019,104
6020,104
6021,104
6022,104
6023,104
6024,104
6025,104
6026,104
6027,104
6028,104
6029,104
6030,104
6031,104
6032,104
6033,104
6034,104
6035,104
6036,104
6037,104
6038,104
6039,104
6040,104
6041,104
6042,105
6043,105
6044,105
6045,105
6046,105
6047,105
6048,105
6049,105
6050,105
6051,105
6052,105
6053,105
6054,105
6055,105
6056,105
6057,105
6058,105
6059,105
6060,105
6061,105
6062,105
6063,105
6064,105
6065,105
6066,105
6067,105
6068,105
6069,105
6070,105
6071,105
6072,105
6073,105
6074,105
6075,105
6076,105
6077,105
6078,105
6079,105
6080,105
6081,105
6082,105
6083,105
6084,105
6085,105
6086,105
6087,105
6088,105
6089,105
6090,105
6091,105
6092,105
6093,105
6094,105
6095,105
6096,105
6097,105
6098,105
6099,105
6100,106
6101,106
6102,106
6103,106
6104,106
6105,106
6106,106
6107,106
6108,106
6109,106
6110,106
6111,106
6112,106
6113,106
6114,106
6115,106
6116,106
6117,106
6118,106
6119,106
6120,106
6121,106
6122,106
6123,106
6124,106
6125,106
6126,106
6127,106
6128,106
6129,106
6130,106
6131,106
6132,106
6133,106
6134,106
6135,106
6136,106
6137,106
6138,106
6139,106
6140,106
6141,106
6142,106
6143,106
6144,106
6145,106
6146,106
6147,106
6148,106
6149,106
6150,106
6151,106
6152,106
6153,106
6154,106
6155,106
6156,106
6157,106
6158,107
6159,107
6160,107
6161,107
6162,107
6163,107
6164,107
6165,107
6166,107
6167,107
6168,107
6169,107
6170,107
6171,107
6172,107
6173,107
6174,107
6175,107
6176,107
6177,107
6178,107
6179,107
6180,107
6181,107
6182,107
6183,107
6184,107
6185,107
6186,107
6187,107
6188,107
6189,107
6190,107
6191,107
6192,107
6193,107
6194,107
6195,107
6196,107
6197,107
6198,107
6199,107
6200,107
6201,107
6202,107
6203,107
6204,107
6205,107
6206,107
6207,107
6208,107
6209,107
6210,107
6211,107
6212,107
6213,107
6214,107
6215,107
6216,108
6217,108
6218,108
6219,108
6220,108
6221,108
6222,108
6223,108
6224,108
6225,108
6226,108
6227,108
6228,108
6229,108
6230,108
6231,108
6232,108
6233,108
6234,108
6235,108
6236,108
6237,108
6238,108
6239,108
6240,108
6241,108
6242,108
6243,108
6244,108
6245,108
6246,108
6247,108
6248,108
6249,108
6250,108
6251,108
6252,108
6253,108
6254,108
6255,108
6256,108
6257,108
6258,108
6259,108
6260,108
6261,108
6262,108
6263,108
6264,108
6265,108
6266,108
6267,108
6268,108
6269,108
6270,108
6271,108
6272,108
6273,108
6274,109
6275,109
6276,109
6277,109
6278,109
6279,109
6280,109
6281,109
6282,109
6283,109
6284,109
6285,109
6286,109
6287,109
6288,109
6289,109
6290,109
6291,109
6292,109
6293,109
6294,109
6295,109
6296,109
6297,109
6298,109
6299,109
6300,109
6301,109
6302,109
6303,109
6304,109
6305,109
6306,109
6307,109
6308,109
6309,109
6310,109
6311,109
6312,109
6313,109
6314,109
6315,109
6316,109
6317,109
6318,109
6319,109
6320,109
6321,109
6322,109
6323,109
6324,109
6325,109
6326,109
6327,109
6328,109
6329,109
6330,109
6331,109
6332,110
6333,110
6334,110
6335,110
6336,110
6337,110
6338,110
6339,110
6340,110
6341,110
6342,110
6343,110
6344,110
6345,110
6346,110
6347,110
6348,110
6349,110
6350,110
6351,110
6352,110
6353,110
6354,110
6355,110
6356,110
6357,110
6358,110
6359,110
6360,110
6361,110
6362,110
6363,110
6364,110
6365,110
6366,110
6367,110
6368,110
6369,110
6370,110
6371,110
6372,110
6373,110
6374,110
6375,110
6376,110
6377,110
6378,110
6379,110
6380,110
6381,110
6382,110
6383,110
6384,110
6385,110
6386,110
6387,110
6388,110
6389,110
6390,111
6391,111
6392,111
6393,111
6394,111
6395,111
6396,111
6397,111
6398,111
6399,111
6400,111
6401,111
6402,111
6403,111
6404,111
6405,111
6406,111
6407,111
6408,111
6409,111
6410,111
6411,111
6412,111
6413,111
6414,111
6415,111
6416,111
6417,111
6418,111
6419,111
6420,111
6421,111
6422,111
6423,111
6424,111
6425,111
6426,111
6427,111
6428,111
6429,111
6430,111
6431,111
6432,111
6433,111
6434,111
6435,111
6436,111
6437,111
6438,111
6439,111
6440,111
6441,111
6442,111
6443,111
6444,111
6445,111
6446,111
6447,111
6448,112
6449,112
6450,112
6451,112
6452,112
6453,112
6454,112
6455,112
6456,112
6457,112
6458,112
6459,112
6460,112
6461,112
6462,112
6463,112
6464,112
6465,112
6466,112
6467,112
6468,112
6469,112
6470,112
6471,112
6472,112
6473,112
6474,112
6475,112
6476,112
6477,112
6478,112
6479,112
6480,112
6481,112
6482,112
6483,112
6484,112
6485,112
6486,112
6487,112
6488,112
6489,112
6490,112
6491,112
6492,112
6493,112
6494,112
6495,112
6496,112
6497,112
6498,112
6499,112
6500,112
6501,112
6502,112
6503,112
6504,112
6505,112
6506,113
6507,113
6508,113
6509,113
6510,113
6511,113
6512,113
6513,113
6514,113
6515,113
6516,113
6517,113
6518,113
6519,113
6520,113
6521,113
6522,113
6523,113
6524,113
6525,113
6526,113
6527,113
6528,113
6529,113
6530,113
6531,113
6532,113
6533,113
6534,113
6535,113
6536,113
6537,113
6538,113
6539,113
6540,113
6541,113
6542,113
6543,113
6544,113
6545,113
6546,113
6547,113
6548,113
6549,113
6550,113
6551,113
6552,113
6553,113
6554,113
6555,113
6556,113
6557,113
6558,113
6559,113
6560,113
6561,113
6562,113
6563,113
6564,114
6565,114
6566,114
6567,114
6568,114
6569,114
6570,114
6571,114
6572,114
6573,114
6574,114
6575,114
6576,114
6577,114
6578,114
6579,114
6580,114
6581,114
6582,114
6583,114
6584,114
6585,114
6586,114
6587,114
6588,114
6589,114
6590,114
6591,114
6592,114
6593,114
6594,114
6595,114
6596,114
6597,114
6598,114
6599,114
6600,114
6601,114
6602,114
6603,114
6604,114
6605,114
6606,114
6607,114
6608,114
6609,114
6610,114
6611,114
6612,114
6613,114
6614,114
6615,114
6616,114
6617,114
6618,114
6619,114
6620,114
6621,114
6622,115
6623,115
6624,115
6625,115
6626,115
6627,115
6628,115
6629,115
6630,115
6631,115
6632,115
6633,115
6634,115
6635,115
6636,115
6637,115
6638,115
6639,115
6640,115
6641,115
6642,115
6643,115
6644,115
6645,115
6646,115
6647,115
6648,115
6649,115
6650,115
6651,115
6652,115
6653,115
6654,115
6655,115
6656,115
6657,115
6658,115
6659,115
6660,115
6661,115
6662,115
6663,115
6664,115
6665,115
6666,115
6667,115
6668,115
6669,115
6670,115
6671,115
6672,115
6673,115
6674,115
6675,115
6676,115
6677,115
6678,115
6679,115
6680,116
6681,116
6682,116
6683,116
6684,116
6685,116
6686,116
6687,116
6688,116
6689,116
6690,116
6691,116
6692,116
6693,116
6694,116
6695,116
6696,116
6697,116
6698,116
6699,116
6700,116
6701,116
6702,116
6703,116
6704,116
6705,116
6706,116
6707,116
6708,116
6709,116
6710,116
6711,116
6712,116
6713,116
6714,116
6715,116
6716,116
6717,116
6718,116
6719,116
6720,116
6721,116
6722,116
6723,116
6724,116
6725,116
6726,116
6727,116
6728,116
6729,116
6730,116
6731,116
6732,116
6733,116
6734,116
6735,116
6736,116
6737,116
6738,117
6739,117
6740,117
6741,117
6742,117
6743,117
6744,117
6745,117
6746,117
6747,117
6748,117
6749,117
6750,117
6751,117
6752,117
6753,117
6754,117
6755,117
6756,117
6757,117
6758,117
6759,117
6760,117
6761,117
6762,117
6763,117
6764,117
6765,117
6766,117
6767,117
6768,117
6769,117
6770,117
6771,117
6772,117
6773,117
6774,117
6775,117
6776,117
6777,117
6778,117
6779,117
6780,117
6781,117
6782,117
6783,117
6784,117
6785,117
6786,117
6787,117
6788,117
6789,117
6790,117
6791,117
6792,117
6793,117
6794,117
6795,117
6796,118
6797,118
6798,118
6799,118
6800,118
6801,118
6802,118
6803,118
6804,118
6805,118
6806,118
6807,118
6808,118
6809,118
6810,118
6811,118
6812,118
6813,118
6814,118
6815,118
6816,118
6817,118
6818,118
6819,118
6820,118
6821,118
6822,118
6823,118
6824,118
6825,118
6826,118
6827,118
6828,118
6829,118
6830,118
6831,118
6832,118
6833,118
6834,118
6835,118
6836,118
6837,118
6838,118
6839,118
6840,118
6841,118
6842,118
6843,118
6844,118
6845,118
6846,118
6847,118
6848,118
6849,118
6850,118
6851,118
6852,118
6853,118
6854,119
6855,119
6856,119
6857,119
6858,119
6859,119
6860,119
6861,119
6862,119
6863,119
6864,119
6865,119
6866,119
6867,119
6868,119
6869,119
6870,119
6871,119
6872,119
6873,119
6874,119
6875,119
6876,119
6877,119
6878,119
6879,119
6880,119
6881,119
6882,119
6883,119
6884,119
6885,119
6886,119
6887,119
6888,119
6889,119
6890,119
6891,119
6892,119
6893,119
6894,119
6895,119
6896,119
6897,119
6898,119
6899,119
6900,119
6901,119
6902,119
6903,119
6904,119
6905,119
6906,119
6907,119
6908,119
6909,119
6910,119
6911,119
