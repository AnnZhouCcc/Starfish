0,0
1,0
2,0
3,0
4,0
5,0
6,0
7,0
8,0
9,0
10,0
11,0
12,0
13,0
14,0
15,0
16,0
17,0
18,0
19,0
20,0
21,0
22,0
23,0
24,0
25,0
26,0
27,0
28,0
29,0
30,0
31,0
32,0
33,0
34,0
35,0
36,0
37,0
38,0
39,0
40,0
41,0
42,0
43,0
44,0
45,0
46,1
47,1
48,1
49,1
50,1
51,1
52,1
53,1
54,1
55,1
56,1
57,1
58,1
59,1
60,1
61,1
62,1
63,1
64,1
65,1
66,1
67,1
68,1
69,1
70,1
71,1
72,1
73,1
74,1
75,1
76,1
77,1
78,1
79,1
80,1
81,1
82,1
83,1
84,1
85,1
86,1
87,1
88,1
89,1
90,1
91,1
92,2
93,2
94,2
95,2
96,2
97,2
98,2
99,2
100,2
101,2
102,2
103,2
104,2
105,2
106,2
107,2
108,2
109,2
110,2
111,2
112,2
113,2
114,2
115,2
116,2
117,2
118,2
119,2
120,2
121,2
122,2
123,2
124,2
125,2
126,2
127,2
128,2
129,2
130,2
131,2
132,2
133,2
134,2
135,2
136,2
137,2
138,3
139,3
140,3
141,3
142,3
143,3
144,3
145,3
146,3
147,3
148,3
149,3
150,3
151,3
152,3
153,3
154,3
155,3
156,3
157,3
158,3
159,3
160,3
161,3
162,3
163,3
164,3
165,3
166,3
167,3
168,3
169,3
170,3
171,3
172,3
173,3
174,3
175,3
176,3
177,3
178,3
179,3
180,3
181,3
182,3
183,3
184,4
185,4
186,4
187,4
188,4
189,4
190,4
191,4
192,4
193,4
194,4
195,4
196,4
197,4
198,4
199,4
200,4
201,4
202,4
203,4
204,4
205,4
206,4
207,4
208,4
209,4
210,4
211,4
212,4
213,4
214,4
215,4
216,4
217,4
218,4
219,4
220,4
221,4
222,4
223,4
224,4
225,4
226,4
227,4
228,4
229,4
230,5
231,5
232,5
233,5
234,5
235,5
236,5
237,5
238,5
239,5
240,5
241,5
242,5
243,5
244,5
245,5
246,5
247,5
248,5
249,5
250,5
251,5
252,5
253,5
254,5
255,5
256,5
257,5
258,5
259,5
260,5
261,5
262,5
263,5
264,5
265,5
266,5
267,5
268,5
269,5
270,5
271,5
272,5
273,5
274,5
275,5
276,6
277,6
278,6
279,6
280,6
281,6
282,6
283,6
284,6
285,6
286,6
287,6
288,6
289,6
290,6
291,6
292,6
293,6
294,6
295,6
296,6
297,6
298,6
299,6
300,6
301,6
302,6
303,6
304,6
305,6
306,6
307,6
308,6
309,6
310,6
311,6
312,6
313,6
314,6
315,6
316,6
317,6
318,6
319,6
320,6
321,6
322,7
323,7
324,7
325,7
326,7
327,7
328,7
329,7
330,7
331,7
332,7
333,7
334,7
335,7
336,7
337,7
338,7
339,7
340,7
341,7
342,7
343,7
344,7
345,7
346,7
347,7
348,7
349,7
350,7
351,7
352,7
353,7
354,7
355,7
356,7
357,7
358,7
359,7
360,7
361,7
362,7
363,7
364,7
365,7
366,7
367,7
368,8
369,8
370,8
371,8
372,8
373,8
374,8
375,8
376,8
377,8
378,8
379,8
380,8
381,8
382,8
383,8
384,8
385,8
386,8
387,8
388,8
389,8
390,8
391,8
392,8
393,8
394,8
395,8
396,8
397,8
398,8
399,8
400,8
401,8
402,8
403,8
404,8
405,8
406,8
407,8
408,8
409,8
410,8
411,8
412,8
413,8
414,9
415,9
416,9
417,9
418,9
419,9
420,9
421,9
422,9
423,9
424,9
425,9
426,9
427,9
428,9
429,9
430,9
431,9
432,9
433,9
434,9
435,9
436,9
437,9
438,9
439,9
440,9
441,9
442,9
443,9
444,9
445,9
446,9
447,9
448,9
449,9
450,9
451,9
452,9
453,9
454,9
455,9
456,9
457,9
458,9
459,9
460,10
461,10
462,10
463,10
464,10
465,10
466,10
467,10
468,10
469,10
470,10
471,10
472,10
473,10
474,10
475,10
476,10
477,10
478,10
479,10
480,10
481,10
482,10
483,10
484,10
485,10
486,10
487,10
488,10
489,10
490,10
491,10
492,10
493,10
494,10
495,10
496,10
497,10
498,10
499,10
500,10
501,10
502,10
503,10
504,10
505,10
506,11
507,11
508,11
509,11
510,11
511,11
512,11
513,11
514,11
515,11
516,11
517,11
518,11
519,11
520,11
521,11
522,11
523,11
524,11
525,11
526,11
527,11
528,11
529,11
530,11
531,11
532,11
533,11
534,11
535,11
536,11
537,11
538,11
539,11
540,11
541,11
542,11
543,11
544,11
545,11
546,11
547,11
548,11
549,11
550,11
551,11
552,12
553,12
554,12
555,12
556,12
557,12
558,12
559,12
560,12
561,12
562,12
563,12
564,12
565,12
566,12
567,12
568,12
569,12
570,12
571,12
572,12
573,12
574,12
575,12
576,12
577,12
578,12
579,12
580,12
581,12
582,12
583,12
584,12
585,12
586,12
587,12
588,12
589,12
590,12
591,12
592,12
593,12
594,12
595,12
596,12
597,12
598,13
599,13
600,13
601,13
602,13
603,13
604,13
605,13
606,13
607,13
608,13
609,13
610,13
611,13
612,13
613,13
614,13
615,13
616,13
617,13
618,13
619,13
620,13
621,13
622,13
623,13
624,13
625,13
626,13
627,13
628,13
629,13
630,13
631,13
632,13
633,13
634,13
635,13
636,13
637,13
638,13
639,13
640,13
641,13
642,13
643,13
644,14
645,14
646,14
647,14
648,14
649,14
650,14
651,14
652,14
653,14
654,14
655,14
656,14
657,14
658,14
659,14
660,14
661,14
662,14
663,14
664,14
665,14
666,14
667,14
668,14
669,14
670,14
671,14
672,14
673,14
674,14
675,14
676,14
677,14
678,14
679,14
680,14
681,14
682,14
683,14
684,14
685,14
686,14
687,14
688,14
689,14
690,15
691,15
692,15
693,15
694,15
695,15
696,15
697,15
698,15
699,15
700,15
701,15
702,15
703,15
704,15
705,15
706,15
707,15
708,15
709,15
710,15
711,15
712,15
713,15
714,15
715,15
716,15
717,15
718,15
719,15
720,15
721,15
722,15
723,15
724,15
725,15
726,15
727,15
728,15
729,15
730,15
731,15
732,15
733,15
734,15
735,15
736,16
737,16
738,16
739,16
740,16
741,16
742,16
743,16
744,16
745,16
746,16
747,16
748,16
749,16
750,16
751,16
752,16
753,16
754,16
755,16
756,16
757,16
758,16
759,16
760,16
761,16
762,16
763,16
764,16
765,16
766,16
767,16
768,16
769,16
770,16
771,16
772,16
773,16
774,16
775,16
776,16
777,16
778,16
779,16
780,16
781,16
782,16
783,16
784,17
785,17
786,17
787,17
788,17
789,17
790,17
791,17
792,17
793,17
794,17
795,17
796,17
797,17
798,17
799,17
800,17
801,17
802,17
803,17
804,17
805,17
806,17
807,17
808,17
809,17
810,17
811,17
812,17
813,17
814,17
815,17
816,17
817,17
818,17
819,17
820,17
821,17
822,17
823,17
824,17
825,17
826,17
827,17
828,17
829,17
830,17
831,17
832,18
833,18
834,18
835,18
836,18
837,18
838,18
839,18
840,18
841,18
842,18
843,18
844,18
845,18
846,18
847,18
848,18
849,18
850,18
851,18
852,18
853,18
854,18
855,18
856,18
857,18
858,18
859,18
860,18
861,18
862,18
863,18
864,18
865,18
866,18
867,18
868,18
869,18
870,18
871,18
872,18
873,18
874,18
875,18
876,18
877,18
878,18
879,18
880,19
881,19
882,19
883,19
884,19
885,19
886,19
887,19
888,19
889,19
890,19
891,19
892,19
893,19
894,19
895,19
896,19
897,19
898,19
899,19
900,19
901,19
902,19
903,19
904,19
905,19
906,19
907,19
908,19
909,19
910,19
911,19
912,19
913,19
914,19
915,19
916,19
917,19
918,19
919,19
920,19
921,19
922,19
923,19
924,19
925,19
926,19
927,19
928,20
929,20
930,20
931,20
932,20
933,20
934,20
935,20
936,20
937,20
938,20
939,20
940,20
941,20
942,20
943,20
944,20
945,20
946,20
947,20
948,20
949,20
950,20
951,20
952,20
953,20
954,20
955,20
956,20
957,20
958,20
959,20
960,20
961,20
962,20
963,20
964,20
965,20
966,20
967,20
968,20
969,20
970,20
971,20
972,20
973,20
974,20
975,20
976,21
977,21
978,21
979,21
980,21
981,21
982,21
983,21
984,21
985,21
986,21
987,21
988,21
989,21
990,21
991,21
992,21
993,21
994,21
995,21
996,21
997,21
998,21
999,21
1000,21
1001,21
1002,21
1003,21
1004,21
1005,21
1006,21
1007,21
1008,21
1009,21
1010,21
1011,21
1012,21
1013,21
1014,21
1015,21
1016,21
1017,21
1018,21
1019,21
1020,21
1021,21
1022,21
1023,21
1024,22
1025,22
1026,22
1027,22
1028,22
1029,22
1030,22
1031,22
1032,22
1033,22
1034,22
1035,22
1036,22
1037,22
1038,22
1039,22
1040,22
1041,22
1042,22
1043,22
1044,22
1045,22
1046,22
1047,22
1048,22
1049,22
1050,22
1051,22
1052,22
1053,22
1054,22
1055,22
1056,22
1057,22
1058,22
1059,22
1060,22
1061,22
1062,22
1063,22
1064,22
1065,22
1066,22
1067,22
1068,22
1069,22
1070,22
1071,22
1072,23
1073,23
1074,23
1075,23
1076,23
1077,23
1078,23
1079,23
1080,23
1081,23
1082,23
1083,23
1084,23
1085,23
1086,23
1087,23
1088,23
1089,23
1090,23
1091,23
1092,23
1093,23
1094,23
1095,23
1096,23
1097,23
1098,23
1099,23
1100,23
1101,23
1102,23
1103,23
1104,23
1105,23
1106,23
1107,23
1108,23
1109,23
1110,23
1111,23
1112,23
1113,23
1114,23
1115,23
1116,23
1117,23
1118,23
1119,23
1120,24
1121,24
1122,24
1123,24
1124,24
1125,24
1126,24
1127,24
1128,24
1129,24
1130,24
1131,24
1132,24
1133,24
1134,24
1135,24
1136,24
1137,24
1138,24
1139,24
1140,24
1141,24
1142,24
1143,24
1144,24
1145,24
1146,24
1147,24
1148,24
1149,24
1150,24
1151,24
1152,24
1153,24
1154,24
1155,24
1156,24
1157,24
1158,24
1159,24
1160,24
1161,24
1162,24
1163,24
1164,24
1165,24
1166,24
1167,24
1168,25
1169,25
1170,25
1171,25
1172,25
1173,25
1174,25
1175,25
1176,25
1177,25
1178,25
1179,25
1180,25
1181,25
1182,25
1183,25
1184,25
1185,25
1186,25
1187,25
1188,25
1189,25
1190,25
1191,25
1192,25
1193,25
1194,25
1195,25
1196,25
1197,25
1198,25
1199,25
1200,25
1201,25
1202,25
1203,25
1204,25
1205,25
1206,25
1207,25
1208,25
1209,25
1210,25
1211,25
1212,25
1213,25
1214,26
1215,26
1216,26
1217,26
1218,26
1219,26
1220,26
1221,26
1222,26
1223,26
1224,26
1225,26
1226,26
1227,26
1228,26
1229,26
1230,26
1231,26
1232,26
1233,26
1234,26
1235,26
1236,26
1237,26
1238,26
1239,26
1240,26
1241,26
1242,26
1243,26
1244,26
1245,26
1246,26
1247,26
1248,26
1249,26
1250,26
1251,26
1252,26
1253,26
1254,26
1255,26
1256,26
1257,26
1258,26
1259,26
1260,27
1261,27
1262,27
1263,27
1264,27
1265,27
1266,27
1267,27
1268,27
1269,27
1270,27
1271,27
1272,27
1273,27
1274,27
1275,27
1276,27
1277,27
1278,27
1279,27
1280,27
1281,27
1282,27
1283,27
1284,27
1285,27
1286,27
1287,27
1288,27
1289,27
1290,27
1291,27
1292,27
1293,27
1294,27
1295,27
1296,27
1297,27
1298,27
1299,27
1300,27
1301,27
1302,27
1303,27
1304,27
1305,27
1306,28
1307,28
1308,28
1309,28
1310,28
1311,28
1312,28
1313,28
1314,28
1315,28
1316,28
1317,28
1318,28
1319,28
1320,28
1321,28
1322,28
1323,28
1324,28
1325,28
1326,28
1327,28
1328,28
1329,28
1330,28
1331,28
1332,28
1333,28
1334,28
1335,28
1336,28
1337,28
1338,28
1339,28
1340,28
1341,28
1342,28
1343,28
1344,28
1345,28
1346,28
1347,28
1348,28
1349,28
1350,28
1351,28
1352,29
1353,29
1354,29
1355,29
1356,29
1357,29
1358,29
1359,29
1360,29
1361,29
1362,29
1363,29
1364,29
1365,29
1366,29
1367,29
1368,29
1369,29
1370,29
1371,29
1372,29
1373,29
1374,29
1375,29
1376,29
1377,29
1378,29
1379,29
1380,29
1381,29
1382,29
1383,29
1384,29
1385,29
1386,29
1387,29
1388,29
1389,29
1390,29
1391,29
1392,29
1393,29
1394,29
1395,29
1396,29
1397,29
1398,30
1399,30
1400,30
1401,30
1402,30
1403,30
1404,30
1405,30
1406,30
1407,30
1408,30
1409,30
1410,30
1411,30
1412,30
1413,30
1414,30
1415,30
1416,30
1417,30
1418,30
1419,30
1420,30
1421,30
1422,30
1423,30
1424,30
1425,30
1426,30
1427,30
1428,30
1429,30
1430,30
1431,30
1432,30
1433,30
1434,30
1435,30
1436,30
1437,30
1438,30
1439,30
1440,30
1441,30
1442,30
1443,30
1444,31
1445,31
1446,31
1447,31
1448,31
1449,31
1450,31
1451,31
1452,31
1453,31
1454,31
1455,31
1456,31
1457,31
1458,31
1459,31
1460,31
1461,31
1462,31
1463,31
1464,31
1465,31
1466,31
1467,31
1468,31
1469,31
1470,31
1471,31
1472,31
1473,31
1474,31
1475,31
1476,31
1477,31
1478,31
1479,31
1480,31
1481,31
1482,31
1483,31
1484,31
1485,31
1486,31
1487,31
1488,31
1489,31
1490,32
1491,32
1492,32
1493,32
1494,32
1495,32
1496,32
1497,32
1498,32
1499,32
1500,32
1501,32
1502,32
1503,32
1504,32
1505,32
1506,32
1507,32
1508,32
1509,32
1510,32
1511,32
1512,32
1513,32
1514,32
1515,32
1516,32
1517,32
1518,32
1519,32
1520,32
1521,32
1522,32
1523,32
1524,32
1525,32
1526,32
1527,32
1528,32
1529,32
1530,32
1531,32
1532,32
1533,32
1534,32
1535,32
1536,33
1537,33
1538,33
1539,33
1540,33
1541,33
1542,33
1543,33
1544,33
1545,33
1546,33
1547,33
1548,33
1549,33
1550,33
1551,33
1552,33
1553,33
1554,33
1555,33
1556,33
1557,33
1558,33
1559,33
1560,33
1561,33
1562,33
1563,33
1564,33
1565,33
1566,33
1567,33
1568,33
1569,33
1570,33
1571,33
1572,33
1573,33
1574,33
1575,33
1576,33
1577,33
1578,33
1579,33
1580,33
1581,33
1582,34
1583,34
1584,34
1585,34
1586,34
1587,34
1588,34
1589,34
1590,34
1591,34
1592,34
1593,34
1594,34
1595,34
1596,34
1597,34
1598,34
1599,34
1600,34
1601,34
1602,34
1603,34
1604,34
1605,34
1606,34
1607,34
1608,34
1609,34
1610,34
1611,34
1612,34
1613,34
1614,34
1615,34
1616,34
1617,34
1618,34
1619,34
1620,34
1621,34
1622,34
1623,34
1624,34
1625,34
1626,34
1627,34
1628,35
1629,35
1630,35
1631,35
1632,35
1633,35
1634,35
1635,35
1636,35
1637,35
1638,35
1639,35
1640,35
1641,35
1642,35
1643,35
1644,35
1645,35
1646,35
1647,35
1648,35
1649,35
1650,35
1651,35
1652,35
1653,35
1654,35
1655,35
1656,35
1657,35
1658,35
1659,35
1660,35
1661,35
1662,35
1663,35
1664,35
1665,35
1666,35
1667,35
1668,35
1669,35
1670,35
1671,35
1672,35
1673,35
1674,36
1675,36
1676,36
1677,36
1678,36
1679,36
1680,36
1681,36
1682,36
1683,36
1684,36
1685,36
1686,36
1687,36
1688,36
1689,36
1690,36
1691,36
1692,36
1693,36
1694,36
1695,36
1696,36
1697,36
1698,36
1699,36
1700,36
1701,36
1702,36
1703,36
1704,36
1705,36
1706,36
1707,36
1708,36
1709,36
1710,36
1711,36
1712,36
1713,36
1714,36
1715,36
1716,36
1717,36
1718,36
1719,36
1720,37
1721,37
1722,37
1723,37
1724,37
1725,37
1726,37
1727,37
1728,37
1729,37
1730,37
1731,37
1732,37
1733,37
1734,37
1735,37
1736,37
1737,37
1738,37
1739,37
1740,37
1741,37
1742,37
1743,37
1744,37
1745,37
1746,37
1747,37
1748,37
1749,37
1750,37
1751,37
1752,37
1753,37
1754,37
1755,37
1756,37
1757,37
1758,37
1759,37
1760,37
1761,37
1762,37
1763,37
1764,37
1765,37
1766,38
1767,38
1768,38
1769,38
1770,38
1771,38
1772,38
1773,38
1774,38
1775,38
1776,38
1777,38
1778,38
1779,38
1780,38
1781,38
1782,38
1783,38
1784,38
1785,38
1786,38
1787,38
1788,38
1789,38
1790,38
1791,38
1792,38
1793,38
1794,38
1795,38
1796,38
1797,38
1798,38
1799,38
1800,38
1801,38
1802,38
1803,38
1804,38
1805,38
1806,38
1807,38
1808,38
1809,38
1810,38
1811,38
1812,39
1813,39
1814,39
1815,39
1816,39
1817,39
1818,39
1819,39
1820,39
1821,39
1822,39
1823,39
1824,39
1825,39
1826,39
1827,39
1828,39
1829,39
1830,39
1831,39
1832,39
1833,39
1834,39
1835,39
1836,39
1837,39
1838,39
1839,39
1840,39
1841,39
1842,39
1843,39
1844,39
1845,39
1846,39
1847,39
1848,39
1849,39
1850,39
1851,39
1852,39
1853,39
1854,39
1855,39
1856,39
1857,39
1858,40
1859,40
1860,40
1861,40
1862,40
1863,40
1864,40
1865,40
1866,40
1867,40
1868,40
1869,40
1870,40
1871,40
1872,40
1873,40
1874,40
1875,40
1876,40
1877,40
1878,40
1879,40
1880,40
1881,40
1882,40
1883,40
1884,40
1885,40
1886,40
1887,40
1888,40
1889,40
1890,40
1891,40
1892,40
1893,40
1894,40
1895,40
1896,40
1897,40
1898,40
1899,40
1900,40
1901,40
1902,40
1903,40
1904,41
1905,41
1906,41
1907,41
1908,41
1909,41
1910,41
1911,41
1912,41
1913,41
1914,41
1915,41
1916,41
1917,41
1918,41
1919,41
1920,41
1921,41
1922,41
1923,41
1924,41
1925,41
1926,41
1927,41
1928,41
1929,41
1930,41
1931,41
1932,41
1933,41
1934,41
1935,41
1936,41
1937,41
1938,41
1939,41
1940,41
1941,41
1942,41
1943,41
1944,41
1945,41
1946,41
1947,41
1948,41
1949,41
1950,41
1951,41
1952,42
1953,42
1954,42
1955,42
1956,42
1957,42
1958,42
1959,42
1960,42
1961,42
1962,42
1963,42
1964,42
1965,42
1966,42
1967,42
1968,42
1969,42
1970,42
1971,42
1972,42
1973,42
1974,42
1975,42
1976,42
1977,42
1978,42
1979,42
1980,42
1981,42
1982,42
1983,42
1984,42
1985,42
1986,42
1987,42
1988,42
1989,42
1990,42
1991,42
1992,42
1993,42
1994,42
1995,42
1996,42
1997,42
1998,42
1999,42
2000,43
2001,43
2002,43
2003,43
2004,43
2005,43
2006,43
2007,43
2008,43
2009,43
2010,43
2011,43
2012,43
2013,43
2014,43
2015,43
2016,43
2017,43
2018,43
2019,43
2020,43
2021,43
2022,43
2023,43
2024,43
2025,43
2026,43
2027,43
2028,43
2029,43
2030,43
2031,43
2032,43
2033,43
2034,43
2035,43
2036,43
2037,43
2038,43
2039,43
2040,43
2041,43
2042,43
2043,43
2044,43
2045,43
2046,43
2047,43
2048,44
2049,44
2050,44
2051,44
2052,44
2053,44
2054,44
2055,44
2056,44
2057,44
2058,44
2059,44
2060,44
2061,44
2062,44
2063,44
2064,44
2065,44
2066,44
2067,44
2068,44
2069,44
2070,44
2071,44
2072,44
2073,44
2074,44
2075,44
2076,44
2077,44
2078,44
2079,44
2080,44
2081,44
2082,44
2083,44
2084,44
2085,44
2086,44
2087,44
2088,44
2089,44
2090,44
2091,44
2092,44
2093,44
2094,44
2095,44
2096,45
2097,45
2098,45
2099,45
2100,45
2101,45
2102,45
2103,45
2104,45
2105,45
2106,45
2107,45
2108,45
2109,45
2110,45
2111,45
2112,45
2113,45
2114,45
2115,45
2116,45
2117,45
2118,45
2119,45
2120,45
2121,45
2122,45
2123,45
2124,45
2125,45
2126,45
2127,45
2128,45
2129,45
2130,45
2131,45
2132,45
2133,45
2134,45
2135,45
2136,45
2137,45
2138,45
2139,45
2140,45
2141,45
2142,45
2143,45
2144,46
2145,46
2146,46
2147,46
2148,46
2149,46
2150,46
2151,46
2152,46
2153,46
2154,46
2155,46
2156,46
2157,46
2158,46
2159,46
2160,46
2161,46
2162,46
2163,46
2164,46
2165,46
2166,46
2167,46
2168,46
2169,46
2170,46
2171,46
2172,46
2173,46
2174,46
2175,46
2176,46
2177,46
2178,46
2179,46
2180,46
2181,46
2182,46
2183,46
2184,46
2185,46
2186,46
2187,46
2188,46
2189,46
2190,46
2191,46
2192,47
2193,47
2194,47
2195,47
2196,47
2197,47
2198,47
2199,47
2200,47
2201,47
2202,47
2203,47
2204,47
2205,47
2206,47
2207,47
2208,47
2209,47
2210,47
2211,47
2212,47
2213,47
2214,47
2215,47
2216,47
2217,47
2218,47
2219,47
2220,47
2221,47
2222,47
2223,47
2224,47
2225,47
2226,47
2227,47
2228,47
2229,47
2230,47
2231,47
2232,47
2233,47
2234,47
2235,47
2236,47
2237,47
2238,47
2239,47
2240,48
2241,48
2242,48
2243,48
2244,48
2245,48
2246,48
2247,48
2248,48
2249,48
2250,48
2251,48
2252,48
2253,48
2254,48
2255,48
2256,48
2257,48
2258,48
2259,48
2260,48
2261,48
2262,48
2263,48
2264,48
2265,48
2266,48
2267,48
2268,48
2269,48
2270,48
2271,48
2272,48
2273,48
2274,48
2275,48
2276,48
2277,48
2278,48
2279,48
2280,48
2281,48
2282,48
2283,48
2284,48
2285,48
2286,48
2287,48
2288,49
2289,49
2290,49
2291,49
2292,49
2293,49
2294,49
2295,49
2296,49
2297,49
2298,49
2299,49
2300,49
2301,49
2302,49
2303,49
2304,49
2305,49
2306,49
2307,49
2308,49
2309,49
2310,49
2311,49
2312,49
2313,49
2314,49
2315,49
2316,49
2317,49
2318,49
2319,49
2320,49
2321,49
2322,49
2323,49
2324,49
2325,49
2326,49
2327,49
2328,49
2329,49
2330,49
2331,49
2332,49
2333,49
2334,49
2335,49
2336,50
2337,50
2338,50
2339,50
2340,50
2341,50
2342,50
2343,50
2344,50
2345,50
2346,50
2347,50
2348,50
2349,50
2350,50
2351,50
2352,50
2353,50
2354,50
2355,50
2356,50
2357,50
2358,50
2359,50
2360,50
2361,50
2362,50
2363,50
2364,50
2365,50
2366,50
2367,50
2368,50
2369,50
2370,50
2371,50
2372,50
2373,50
2374,50
2375,50
2376,50
2377,50
2378,50
2379,50
2380,50
2381,50
2382,51
2383,51
2384,51
2385,51
2386,51
2387,51
2388,51
2389,51
2390,51
2391,51
2392,51
2393,51
2394,51
2395,51
2396,51
2397,51
2398,51
2399,51
2400,51
2401,51
2402,51
2403,51
2404,51
2405,51
2406,51
2407,51
2408,51
2409,51
2410,51
2411,51
2412,51
2413,51
2414,51
2415,51
2416,51
2417,51
2418,51
2419,51
2420,51
2421,51
2422,51
2423,51
2424,51
2425,51
2426,51
2427,51
2428,52
2429,52
2430,52
2431,52
2432,52
2433,52
2434,52
2435,52
2436,52
2437,52
2438,52
2439,52
2440,52
2441,52
2442,52
2443,52
2444,52
2445,52
2446,52
2447,52
2448,52
2449,52
2450,52
2451,52
2452,52
2453,52
2454,52
2455,52
2456,52
2457,52
2458,52
2459,52
2460,52
2461,52
2462,52
2463,52
2464,52
2465,52
2466,52
2467,52
2468,52
2469,52
2470,52
2471,52
2472,52
2473,52
2474,53
2475,53
2476,53
2477,53
2478,53
2479,53
2480,53
2481,53
2482,53
2483,53
2484,53
2485,53
2486,53
2487,53
2488,53
2489,53
2490,53
2491,53
2492,53
2493,53
2494,53
2495,53
2496,53
2497,53
2498,53
2499,53
2500,53
2501,53
2502,53
2503,53
2504,53
2505,53
2506,53
2507,53
2508,53
2509,53
2510,53
2511,53
2512,53
2513,53
2514,53
2515,53
2516,53
2517,53
2518,53
2519,53
2520,54
2521,54
2522,54
2523,54
2524,54
2525,54
2526,54
2527,54
2528,54
2529,54
2530,54
2531,54
2532,54
2533,54
2534,54
2535,54
2536,54
2537,54
2538,54
2539,54
2540,54
2541,54
2542,54
2543,54
2544,54
2545,54
2546,54
2547,54
2548,54
2549,54
2550,54
2551,54
2552,54
2553,54
2554,54
2555,54
2556,54
2557,54
2558,54
2559,54
2560,54
2561,54
2562,54
2563,54
2564,54
2565,54
2566,55
2567,55
2568,55
2569,55
2570,55
2571,55
2572,55
2573,55
2574,55
2575,55
2576,55
2577,55
2578,55
2579,55
2580,55
2581,55
2582,55
2583,55
2584,55
2585,55
2586,55
2587,55
2588,55
2589,55
2590,55
2591,55
2592,55
2593,55
2594,55
2595,55
2596,55
2597,55
2598,55
2599,55
2600,55
2601,55
2602,55
2603,55
2604,55
2605,55
2606,55
2607,55
2608,55
2609,55
2610,55
2611,55
2612,56
2613,56
2614,56
2615,56
2616,56
2617,56
2618,56
2619,56
2620,56
2621,56
2622,56
2623,56
2624,56
2625,56
2626,56
2627,56
2628,56
2629,56
2630,56
2631,56
2632,56
2633,56
2634,56
2635,56
2636,56
2637,56
2638,56
2639,56
2640,56
2641,56
2642,56
2643,56
2644,56
2645,56
2646,56
2647,56
2648,56
2649,56
2650,56
2651,56
2652,56
2653,56
2654,56
2655,56
2656,56
2657,56
2658,57
2659,57
2660,57
2661,57
2662,57
2663,57
2664,57
2665,57
2666,57
2667,57
2668,57
2669,57
2670,57
2671,57
2672,57
2673,57
2674,57
2675,57
2676,57
2677,57
2678,57
2679,57
2680,57
2681,57
2682,57
2683,57
2684,57
2685,57
2686,57
2687,57
2688,57
2689,57
2690,57
2691,57
2692,57
2693,57
2694,57
2695,57
2696,57
2697,57
2698,57
2699,57
2700,57
2701,57
2702,57
2703,57
2704,58
2705,58
2706,58
2707,58
2708,58
2709,58
2710,58
2711,58
2712,58
2713,58
2714,58
2715,58
2716,58
2717,58
2718,58
2719,58
2720,58
2721,58
2722,58
2723,58
2724,58
2725,58
2726,58
2727,58
2728,58
2729,58
2730,58
2731,58
2732,58
2733,58
2734,58
2735,58
2736,58
2737,58
2738,58
2739,58
2740,58
2741,58
2742,58
2743,58
2744,58
2745,58
2746,58
2747,58
2748,58
2749,58
2750,59
2751,59
2752,59
2753,59
2754,59
2755,59
2756,59
2757,59
2758,59
2759,59
2760,59
2761,59
2762,59
2763,59
2764,59
2765,59
2766,59
2767,59
2768,59
2769,59
2770,59
2771,59
2772,59
2773,59
2774,59
2775,59
2776,59
2777,59
2778,59
2779,59
2780,59
2781,59
2782,59
2783,59
2784,59
2785,59
2786,59
2787,59
2788,59
2789,59
2790,59
2791,59
2792,59
2793,59
2794,59
2795,59
2796,60
2797,60
2798,60
2799,60
2800,60
2801,60
2802,60
2803,60
2804,60
2805,60
2806,60
2807,60
2808,60
2809,60
2810,60
2811,60
2812,60
2813,60
2814,60
2815,60
2816,60
2817,60
2818,60
2819,60
2820,60
2821,60
2822,60
2823,60
2824,60
2825,60
2826,60
2827,60
2828,60
2829,60
2830,60
2831,60
2832,60
2833,60
2834,60
2835,60
2836,60
2837,60
2838,60
2839,60
2840,60
2841,60
2842,61
2843,61
2844,61
2845,61
2846,61
2847,61
2848,61
2849,61
2850,61
2851,61
2852,61
2853,61
2854,61
2855,61
2856,61
2857,61
2858,61
2859,61
2860,61
2861,61
2862,61
2863,61
2864,61
2865,61
2866,61
2867,61
2868,61
2869,61
2870,61
2871,61
2872,61
2873,61
2874,61
2875,61
2876,61
2877,61
2878,61
2879,61
2880,61
2881,61
2882,61
2883,61
2884,61
2885,61
2886,61
2887,61
2888,62
2889,62
2890,62
2891,62
2892,62
2893,62
2894,62
2895,62
2896,62
2897,62
2898,62
2899,62
2900,62
2901,62
2902,62
2903,62
2904,62
2905,62
2906,62
2907,62
2908,62
2909,62
2910,62
2911,62
2912,62
2913,62
2914,62
2915,62
2916,62
2917,62
2918,62
2919,62
2920,62
2921,62
2922,62
2923,62
2924,62
2925,62
2926,62
2927,62
2928,62
2929,62
2930,62
2931,62
2932,62
2933,62
2934,63
2935,63
2936,63
2937,63
2938,63
2939,63
2940,63
2941,63
2942,63
2943,63
2944,63
2945,63
2946,63
2947,63
2948,63
2949,63
2950,63
2951,63
2952,63
2953,63
2954,63
2955,63
2956,63
2957,63
2958,63
2959,63
2960,63
2961,63
2962,63
2963,63
2964,63
2965,63
2966,63
2967,63
2968,63
2969,63
2970,63
2971,63
2972,63
2973,63
2974,63
2975,63
2976,63
2977,63
2978,63
2979,63
2980,64
2981,64
2982,64
2983,64
2984,64
2985,64
2986,64
2987,64
2988,64
2989,64
2990,64
2991,64
2992,64
2993,64
2994,64
2995,64
2996,64
2997,64
2998,64
2999,64
3000,64
3001,64
3002,64
3003,64
3004,64
3005,64
3006,64
3007,64
3008,64
3009,64
3010,64
3011,64
3012,64
3013,64
3014,64
3015,64
3016,64
3017,64
3018,64
3019,64
3020,64
3021,64
3022,64
3023,64
3024,64
3025,64
3026,65
3027,65
3028,65
3029,65
3030,65
3031,65
3032,65
3033,65
3034,65
3035,65
3036,65
3037,65
3038,65
3039,65
3040,65
3041,65
3042,65
3043,65
3044,65
3045,65
3046,65
3047,65
3048,65
3049,65
3050,65
3051,65
3052,65
3053,65
3054,65
3055,65
3056,65
3057,65
3058,65
3059,65
3060,65
3061,65
3062,65
3063,65
3064,65
3065,65
3066,65
3067,65
3068,65
3069,65
3070,65
3071,65
3072,66
3073,66
3074,66
3075,66
3076,66
3077,66
3078,66
3079,66
3080,66
3081,66
3082,66
3083,66
3084,66
3085,66
3086,66
3087,66
3088,66
3089,66
3090,66
3091,66
3092,66
3093,66
3094,66
3095,66
3096,66
3097,66
3098,66
3099,66
3100,66
3101,66
3102,66
3103,66
3104,66
3105,66
3106,66
3107,66
3108,66
3109,66
3110,66
3111,66
3112,66
3113,66
3114,66
3115,66
3116,66
3117,66
3118,66
3119,66
3120,67
3121,67
3122,67
3123,67
3124,67
3125,67
3126,67
3127,67
3128,67
3129,67
3130,67
3131,67
3132,67
3133,67
3134,67
3135,67
3136,67
3137,67
3138,67
3139,67
3140,67
3141,67
3142,67
3143,67
3144,67
3145,67
3146,67
3147,67
3148,67
3149,67
3150,67
3151,67
3152,67
3153,67
3154,67
3155,67
3156,67
3157,67
3158,67
3159,67
3160,67
3161,67
3162,67
3163,67
3164,67
3165,67
3166,67
3167,67
3168,68
3169,68
3170,68
3171,68
3172,68
3173,68
3174,68
3175,68
3176,68
3177,68
3178,68
3179,68
3180,68
3181,68
3182,68
3183,68
3184,68
3185,68
3186,68
3187,68
3188,68
3189,68
3190,68
3191,68
3192,68
3193,68
3194,68
3195,68
3196,68
3197,68
3198,68
3199,68
3200,68
3201,68
3202,68
3203,68
3204,68
3205,68
3206,68
3207,68
3208,68
3209,68
3210,68
3211,68
3212,68
3213,68
3214,68
3215,68
3216,69
3217,69
3218,69
3219,69
3220,69
3221,69
3222,69
3223,69
3224,69
3225,69
3226,69
3227,69
3228,69
3229,69
3230,69
3231,69
3232,69
3233,69
3234,69
3235,69
3236,69
3237,69
3238,69
3239,69
3240,69
3241,69
3242,69
3243,69
3244,69
3245,69
3246,69
3247,69
3248,69
3249,69
3250,69
3251,69
3252,69
3253,69
3254,69
3255,69
3256,69
3257,69
3258,69
3259,69
3260,69
3261,69
3262,69
3263,69
3264,70
3265,70
3266,70
3267,70
3268,70
3269,70
3270,70
3271,70
3272,70
3273,70
3274,70
3275,70
3276,70
3277,70
3278,70
3279,70
3280,70
3281,70
3282,70
3283,70
3284,70
3285,70
3286,70
3287,70
3288,70
3289,70
3290,70
3291,70
3292,70
3293,70
3294,70
3295,70
3296,70
3297,70
3298,70
3299,70
3300,70
3301,70
3302,70
3303,70
3304,70
3305,70
3306,70
3307,70
3308,70
3309,70
3310,70
3311,70
3312,71
3313,71
3314,71
3315,71
3316,71
3317,71
3318,71
3319,71
3320,71
3321,71
3322,71
3323,71
3324,71
3325,71
3326,71
3327,71
3328,71
3329,71
3330,71
3331,71
3332,71
3333,71
3334,71
3335,71
3336,71
3337,71
3338,71
3339,71
3340,71
3341,71
3342,71
3343,71
3344,71
3345,71
3346,71
3347,71
3348,71
3349,71
3350,71
3351,71
3352,71
3353,71
3354,71
3355,71
3356,71
3357,71
3358,71
3359,71
3360,72
3361,72
3362,72
3363,72
3364,72
3365,72
3366,72
3367,72
3368,72
3369,72
3370,72
3371,72
3372,72
3373,72
3374,72
3375,72
3376,72
3377,72
3378,72
3379,72
3380,72
3381,72
3382,72
3383,72
3384,72
3385,72
3386,72
3387,72
3388,72
3389,72
3390,72
3391,72
3392,72
3393,72
3394,72
3395,72
3396,72
3397,72
3398,72
3399,72
3400,72
3401,72
3402,72
3403,72
3404,72
3405,72
3406,72
3407,72
3408,73
3409,73
3410,73
3411,73
3412,73
3413,73
3414,73
3415,73
3416,73
3417,73
3418,73
3419,73
3420,73
3421,73
3422,73
3423,73
3424,73
3425,73
3426,73
3427,73
3428,73
3429,73
3430,73
3431,73
3432,73
3433,73
3434,73
3435,73
3436,73
3437,73
3438,73
3439,73
3440,73
3441,73
3442,73
3443,73
3444,73
3445,73
3446,73
3447,73
3448,73
3449,73
3450,73
3451,73
3452,73
3453,73
3454,73
3455,73
3456,74
3457,74
3458,74
3459,74
3460,74
3461,74
3462,74
3463,74
3464,74
3465,74
3466,74
3467,74
3468,74
3469,74
3470,74
3471,74
3472,74
3473,74
3474,74
3475,74
3476,74
3477,74
3478,74
3479,74
3480,74
3481,74
3482,74
3483,74
3484,74
3485,74
3486,74
3487,74
3488,74
3489,74
3490,74
3491,74
3492,74
3493,74
3494,74
3495,74
3496,74
3497,74
3498,74
3499,74
3500,74
3501,74
3502,74
3503,74
3504,75
3505,75
3506,75
3507,75
3508,75
3509,75
3510,75
3511,75
3512,75
3513,75
3514,75
3515,75
3516,75
3517,75
3518,75
3519,75
3520,75
3521,75
3522,75
3523,75
3524,75
3525,75
3526,75
3527,75
3528,75
3529,75
3530,75
3531,75
3532,75
3533,75
3534,75
3535,75
3536,75
3537,75
3538,75
3539,75
3540,75
3541,75
3542,75
3543,75
3544,75
3545,75
3546,75
3547,75
3548,75
3549,75
3550,76
3551,76
3552,76
3553,76
3554,76
3555,76
3556,76
3557,76
3558,76
3559,76
3560,76
3561,76
3562,76
3563,76
3564,76
3565,76
3566,76
3567,76
3568,76
3569,76
3570,76
3571,76
3572,76
3573,76
3574,76
3575,76
3576,76
3577,76
3578,76
3579,76
3580,76
3581,76
3582,76
3583,76
3584,76
3585,76
3586,76
3587,76
3588,76
3589,76
3590,76
3591,76
3592,76
3593,76
3594,76
3595,76
3596,77
3597,77
3598,77
3599,77
3600,77
3601,77
3602,77
3603,77
3604,77
3605,77
3606,77
3607,77
3608,77
3609,77
3610,77
3611,77
3612,77
3613,77
3614,77
3615,77
3616,77
3617,77
3618,77
3619,77
3620,77
3621,77
3622,77
3623,77
3624,77
3625,77
3626,77
3627,77
3628,77
3629,77
3630,77
3631,77
3632,77
3633,77
3634,77
3635,77
3636,77
3637,77
3638,77
3639,77
3640,77
3641,77
3642,78
3643,78
3644,78
3645,78
3646,78
3647,78
3648,78
3649,78
3650,78
3651,78
3652,78
3653,78
3654,78
3655,78
3656,78
3657,78
3658,78
3659,78
3660,78
3661,78
3662,78
3663,78
3664,78
3665,78
3666,78
3667,78
3668,78
3669,78
3670,78
3671,78
3672,78
3673,78
3674,78
3675,78
3676,78
3677,78
3678,78
3679,78
3680,78
3681,78
3682,78
3683,78
3684,78
3685,78
3686,78
3687,78
3688,79
3689,79
3690,79
3691,79
3692,79
3693,79
3694,79
3695,79
3696,79
3697,79
3698,79
3699,79
3700,79
3701,79
3702,79
3703,79
3704,79
3705,79
3706,79
3707,79
3708,79
3709,79
3710,79
3711,79
3712,79
3713,79
3714,79
3715,79
3716,79
3717,79
3718,79
3719,79
3720,79
3721,79
3722,79
3723,79
3724,79
3725,79
3726,79
3727,79
3728,79
3729,79
3730,79
3731,79
3732,79
3733,79
3734,80
3735,80
3736,80
3737,80
3738,80
3739,80
3740,80
3741,80
3742,80
3743,80
3744,80
3745,80
3746,80
3747,80
3748,80
3749,80
3750,80
3751,80
3752,80
3753,80
3754,80
3755,80
3756,80
3757,80
3758,80
3759,80
3760,80
3761,80
3762,80
3763,80
3764,80
3765,80
3766,80
3767,80
3768,80
3769,80
3770,80
3771,80
3772,80
3773,80
3774,80
3775,80
3776,80
3777,80
3778,80
3779,80
3780,81
3781,81
3782,81
3783,81
3784,81
3785,81
3786,81
3787,81
3788,81
3789,81
3790,81
3791,81
3792,81
3793,81
3794,81
3795,81
3796,81
3797,81
3798,81
3799,81
3800,81
3801,81
3802,81
3803,81
3804,81
3805,81
3806,81
3807,81
3808,81
3809,81
3810,81
3811,81
3812,81
3813,81
3814,81
3815,81
3816,81
3817,81
3818,81
3819,81
3820,81
3821,81
3822,81
3823,81
3824,81
3825,81
3826,82
3827,82
3828,82
3829,82
3830,82
3831,82
3832,82
3833,82
3834,82
3835,82
3836,82
3837,82
3838,82
3839,82
3840,82
3841,82
3842,82
3843,82
3844,82
3845,82
3846,82
3847,82
3848,82
3849,82
3850,82
3851,82
3852,82
3853,82
3854,82
3855,82
3856,82
3857,82
3858,82
3859,82
3860,82
3861,82
3862,82
3863,82
3864,82
3865,82
3866,82
3867,82
3868,82
3869,82
3870,82
3871,82
3872,83
3873,83
3874,83
3875,83
3876,83
3877,83
3878,83
3879,83
3880,83
3881,83
3882,83
3883,83
3884,83
3885,83
3886,83
3887,83
3888,83
3889,83
3890,83
3891,83
3892,83
3893,83
3894,83
3895,83
3896,83
3897,83
3898,83
3899,83
3900,83
3901,83
3902,83
3903,83
3904,83
3905,83
3906,83
3907,83
3908,83
3909,83
3910,83
3911,83
3912,83
3913,83
3914,83
3915,83
3916,83
3917,83
3918,84
3919,84
3920,84
3921,84
3922,84
3923,84
3924,84
3925,84
3926,84
3927,84
3928,84
3929,84
3930,84
3931,84
3932,84
3933,84
3934,84
3935,84
3936,84
3937,84
3938,84
3939,84
3940,84
3941,84
3942,84
3943,84
3944,84
3945,84
3946,84
3947,84
3948,84
3949,84
3950,84
3951,84
3952,84
3953,84
3954,84
3955,84
3956,84
3957,84
3958,84
3959,84
3960,84
3961,84
3962,84
3963,84
3964,85
3965,85
3966,85
3967,85
3968,85
3969,85
3970,85
3971,85
3972,85
3973,85
3974,85
3975,85
3976,85
3977,85
3978,85
3979,85
3980,85
3981,85
3982,85
3983,85
3984,85
3985,85
3986,85
3987,85
3988,85
3989,85
3990,85
3991,85
3992,85
3993,85
3994,85
3995,85
3996,85
3997,85
3998,85
3999,85
4000,85
4001,85
4002,85
4003,85
4004,85
4005,85
4006,85
4007,85
4008,85
4009,85
4010,86
4011,86
4012,86
4013,86
4014,86
4015,86
4016,86
4017,86
4018,86
4019,86
4020,86
4021,86
4022,86
4023,86
4024,86
4025,86
4026,86
4027,86
4028,86
4029,86
4030,86
4031,86
4032,86
4033,86
4034,86
4035,86
4036,86
4037,86
4038,86
4039,86
4040,86
4041,86
4042,86
4043,86
4044,86
4045,86
4046,86
4047,86
4048,86
4049,86
4050,86
4051,86
4052,86
4053,86
4054,86
4055,86
4056,87
4057,87
4058,87
4059,87
4060,87
4061,87
4062,87
4063,87
4064,87
4065,87
4066,87
4067,87
4068,87
4069,87
4070,87
4071,87
4072,87
4073,87
4074,87
4075,87
4076,87
4077,87
4078,87
4079,87
4080,87
4081,87
4082,87
4083,87
4084,87
4085,87
4086,87
4087,87
4088,87
4089,87
4090,87
4091,87
4092,87
4093,87
4094,87
4095,87
4096,87
4097,87
4098,87
4099,87
4100,87
4101,87
4102,88
4103,88
4104,88
4105,88
4106,88
4107,88
4108,88
4109,88
4110,88
4111,88
4112,88
4113,88
4114,88
4115,88
4116,88
4117,88
4118,88
4119,88
4120,88
4121,88
4122,88
4123,88
4124,88
4125,88
4126,88
4127,88
4128,88
4129,88
4130,88
4131,88
4132,88
4133,88
4134,88
4135,88
4136,88
4137,88
4138,88
4139,88
4140,88
4141,88
4142,88
4143,88
4144,88
4145,88
4146,88
4147,88
4148,89
4149,89
4150,89
4151,89
4152,89
4153,89
4154,89
4155,89
4156,89
4157,89
4158,89
4159,89
4160,89
4161,89
4162,89
4163,89
4164,89
4165,89
4166,89
4167,89
4168,89
4169,89
4170,89
4171,89
4172,89
4173,89
4174,89
4175,89
4176,89
4177,89
4178,89
4179,89
4180,89
4181,89
4182,89
4183,89
4184,89
4185,89
4186,89
4187,89
4188,89
4189,89
4190,89
4191,89
4192,89
4193,89
4194,90
4195,90
4196,90
4197,90
4198,90
4199,90
4200,90
4201,90
4202,90
4203,90
4204,90
4205,90
4206,90
4207,90
4208,90
4209,90
4210,90
4211,90
4212,90
4213,90
4214,90
4215,90
4216,90
4217,90
4218,90
4219,90
4220,90
4221,90
4222,90
4223,90
4224,90
4225,90
4226,90
4227,90
4228,90
4229,90
4230,90
4231,90
4232,90
4233,90
4234,90
4235,90
4236,90
4237,90
4238,90
4239,90
4240,91
4241,91
4242,91
4243,91
4244,91
4245,91
4246,91
4247,91
4248,91
4249,91
4250,91
4251,91
4252,91
4253,91
4254,91
4255,91
4256,91
4257,91
4258,91
4259,91
4260,91
4261,91
4262,91
4263,91
4264,91
4265,91
4266,91
4267,91
4268,91
4269,91
4270,91
4271,91
4272,91
4273,91
4274,91
4275,91
4276,91
4277,91
4278,91
4279,91
4280,91
4281,91
4282,91
4283,91
4284,91
4285,91
4286,91
4287,91
4288,92
4289,92
4290,92
4291,92
4292,92
4293,92
4294,92
4295,92
4296,92
4297,92
4298,92
4299,92
4300,92
4301,92
4302,92
4303,92
4304,92
4305,92
4306,92
4307,92
4308,92
4309,92
4310,92
4311,92
4312,92
4313,92
4314,92
4315,92
4316,92
4317,92
4318,92
4319,92
4320,92
4321,92
4322,92
4323,92
4324,92
4325,92
4326,92
4327,92
4328,92
4329,92
4330,92
4331,92
4332,92
4333,92
4334,92
4335,92
4336,93
4337,93
4338,93
4339,93
4340,93
4341,93
4342,93
4343,93
4344,93
4345,93
4346,93
4347,93
4348,93
4349,93
4350,93
4351,93
4352,93
4353,93
4354,93
4355,93
4356,93
4357,93
4358,93
4359,93
4360,93
4361,93
4362,93
4363,93
4364,93
4365,93
4366,93
4367,93
4368,93
4369,93
4370,93
4371,93
4372,93
4373,93
4374,93
4375,93
4376,93
4377,93
4378,93
4379,93
4380,93
4381,93
4382,93
4383,93
4384,94
4385,94
4386,94
4387,94
4388,94
4389,94
4390,94
4391,94
4392,94
4393,94
4394,94
4395,94
4396,94
4397,94
4398,94
4399,94
4400,94
4401,94
4402,94
4403,94
4404,94
4405,94
4406,94
4407,94
4408,94
4409,94
4410,94
4411,94
4412,94
4413,94
4414,94
4415,94
4416,94
4417,94
4418,94
4419,94
4420,94
4421,94
4422,94
4423,94
4424,94
4425,94
4426,94
4427,94
4428,94
4429,94
4430,94
4431,94
4432,95
4433,95
4434,95
4435,95
4436,95
4437,95
4438,95
4439,95
4440,95
4441,95
4442,95
4443,95
4444,95
4445,95
4446,95
4447,95
4448,95
4449,95
4450,95
4451,95
4452,95
4453,95
4454,95
4455,95
4456,95
4457,95
4458,95
4459,95
4460,95
4461,95
4462,95
4463,95
4464,95
4465,95
4466,95
4467,95
4468,95
4469,95
4470,95
4471,95
4472,95
4473,95
4474,95
4475,95
4476,95
4477,95
4478,95
4479,95
4480,96
4481,96
4482,96
4483,96
4484,96
4485,96
4486,96
4487,96
4488,96
4489,96
4490,96
4491,96
4492,96
4493,96
4494,96
4495,96
4496,96
4497,96
4498,96
4499,96
4500,96
4501,96
4502,96
4503,96
4504,96
4505,96
4506,96
4507,96
4508,96
4509,96
4510,96
4511,96
4512,96
4513,96
4514,96
4515,96
4516,96
4517,96
4518,96
4519,96
4520,96
4521,96
4522,96
4523,96
4524,96
4525,96
4526,96
4527,96
4528,97
4529,97
4530,97
4531,97
4532,97
4533,97
4534,97
4535,97
4536,97
4537,97
4538,97
4539,97
4540,97
4541,97
4542,97
4543,97
4544,97
4545,97
4546,97
4547,97
4548,97
4549,97
4550,97
4551,97
4552,97
4553,97
4554,97
4555,97
4556,97
4557,97
4558,97
4559,97
4560,97
4561,97
4562,97
4563,97
4564,97
4565,97
4566,97
4567,97
4568,97
4569,97
4570,97
4571,97
4572,97
4573,97
4574,97
4575,97
4576,98
4577,98
4578,98
4579,98
4580,98
4581,98
4582,98
4583,98
4584,98
4585,98
4586,98
4587,98
4588,98
4589,98
4590,98
4591,98
4592,98
4593,98
4594,98
4595,98
4596,98
4597,98
4598,98
4599,98
4600,98
4601,98
4602,98
4603,98
4604,98
4605,98
4606,98
4607,98
4608,98
4609,98
4610,98
4611,98
4612,98
4613,98
4614,98
4615,98
4616,98
4617,98
4618,98
4619,98
4620,98
4621,98
4622,98
4623,98
4624,99
4625,99
4626,99
4627,99
4628,99
4629,99
4630,99
4631,99
4632,99
4633,99
4634,99
4635,99
4636,99
4637,99
4638,99
4639,99
4640,99
4641,99
4642,99
4643,99
4644,99
4645,99
4646,99
4647,99
4648,99
4649,99
4650,99
4651,99
4652,99
4653,99
4654,99
4655,99
4656,99
4657,99
4658,99
4659,99
4660,99
4661,99
4662,99
4663,99
4664,99
4665,99
4666,99
4667,99
4668,99
4669,99
4670,99
4671,99
