0,0
1,0
2,0
3,0
4,0
5,0
6,0
7,0
8,0
9,0
10,0
11,0
12,0
13,0
14,0
15,0
16,0
17,0
18,0
19,0
20,0
21,0
22,0
23,0
24,0
25,0
26,0
27,0
28,0
29,0
30,0
31,0
32,0
33,0
34,0
35,0
36,0
37,0
38,0
39,0
40,0
41,0
42,0
43,0
44,0
45,0
46,0
47,0
48,1
49,1
50,1
51,1
52,1
53,1
54,1
55,1
56,1
57,1
58,1
59,1
60,1
61,1
62,1
63,1
64,1
65,1
66,1
67,1
68,1
69,1
70,1
71,1
72,1
73,1
74,1
75,1
76,1
77,1
78,1
79,1
80,1
81,1
82,1
83,1
84,1
85,1
86,1
87,1
88,1
89,1
90,1
91,1
92,1
93,1
94,1
95,1
96,2
97,2
98,2
99,2
100,2
101,2
102,2
103,2
104,2
105,2
106,2
107,2
108,2
109,2
110,2
111,2
112,2
113,2
114,2
115,2
116,2
117,2
118,2
119,2
120,2
121,2
122,2
123,2
124,2
125,2
126,2
127,2
128,2
129,2
130,2
131,2
132,2
133,2
134,2
135,2
136,2
137,2
138,2
139,2
140,2
141,2
142,2
143,2
144,3
145,3
146,3
147,3
148,3
149,3
150,3
151,3
152,3
153,3
154,3
155,3
156,3
157,3
158,3
159,3
160,3
161,3
162,3
163,3
164,3
165,3
166,3
167,3
168,3
169,3
170,3
171,3
172,3
173,3
174,3
175,3
176,3
177,3
178,3
179,3
180,3
181,3
182,3
183,3
184,3
185,3
186,3
187,3
188,3
189,3
190,3
191,3
192,4
193,4
194,4
195,4
196,4
197,4
198,4
199,4
200,4
201,4
202,4
203,4
204,4
205,4
206,4
207,4
208,4
209,4
210,4
211,4
212,4
213,4
214,4
215,4
216,4
217,4
218,4
219,4
220,4
221,4
222,4
223,4
224,4
225,4
226,4
227,4
228,4
229,4
230,4
231,4
232,4
233,4
234,4
235,4
236,4
237,4
238,4
239,4
240,5
241,5
242,5
243,5
244,5
245,5
246,5
247,5
248,5
249,5
250,5
251,5
252,5
253,5
254,5
255,5
256,5
257,5
258,5
259,5
260,5
261,5
262,5
263,5
264,5
265,5
266,5
267,5
268,5
269,5
270,5
271,5
272,5
273,5
274,5
275,5
276,5
277,5
278,5
279,5
280,5
281,5
282,5
283,5
284,5
285,5
286,5
287,5
288,6
289,6
290,6
291,6
292,6
293,6
294,6
295,6
296,6
297,6
298,6
299,6
300,6
301,6
302,6
303,6
304,6
305,6
306,6
307,6
308,6
309,6
310,6
311,6
312,6
313,6
314,6
315,6
316,6
317,6
318,6
319,6
320,6
321,6
322,6
323,6
324,6
325,6
326,6
327,6
328,6
329,6
330,6
331,6
332,6
333,6
334,6
335,6
336,7
337,7
338,7
339,7
340,7
341,7
342,7
343,7
344,7
345,7
346,7
347,7
348,7
349,7
350,7
351,7
352,7
353,7
354,7
355,7
356,7
357,7
358,7
359,7
360,7
361,7
362,7
363,7
364,7
365,7
366,7
367,7
368,7
369,7
370,7
371,7
372,7
373,7
374,7
375,7
376,7
377,7
378,7
379,7
380,7
381,7
382,7
383,7
384,8
385,8
386,8
387,8
388,8
389,8
390,8
391,8
392,8
393,8
394,8
395,8
396,8
397,8
398,8
399,8
400,8
401,8
402,8
403,8
404,8
405,8
406,8
407,8
408,8
409,8
410,8
411,8
412,8
413,8
414,8
415,8
416,8
417,8
418,8
419,8
420,8
421,8
422,8
423,8
424,8
425,8
426,8
427,8
428,8
429,8
430,8
431,8
432,9
433,9
434,9
435,9
436,9
437,9
438,9
439,9
440,9
441,9
442,9
443,9
444,9
445,9
446,9
447,9
448,9
449,9
450,9
451,9
452,9
453,9
454,9
455,9
456,9
457,9
458,9
459,9
460,9
461,9
462,9
463,9
464,9
465,9
466,9
467,9
468,9
469,9
470,9
471,9
472,9
473,9
474,9
475,9
476,9
477,9
478,9
479,9
480,10
481,10
482,10
483,10
484,10
485,10
486,10
487,10
488,10
489,10
490,10
491,10
492,10
493,10
494,10
495,10
496,10
497,10
498,10
499,10
500,10
501,10
502,10
503,10
504,10
505,10
506,10
507,10
508,10
509,10
510,10
511,10
512,10
513,10
514,10
515,10
516,10
517,10
518,10
519,10
520,10
521,10
522,10
523,10
524,10
525,10
526,10
527,10
528,11
529,11
530,11
531,11
532,11
533,11
534,11
535,11
536,11
537,11
538,11
539,11
540,11
541,11
542,11
543,11
544,11
545,11
546,11
547,11
548,11
549,11
550,11
551,11
552,11
553,11
554,11
555,11
556,11
557,11
558,11
559,11
560,11
561,11
562,11
563,11
564,11
565,11
566,11
567,11
568,11
569,11
570,11
571,11
572,11
573,11
574,11
575,11
576,12
577,12
578,12
579,12
580,12
581,12
582,12
583,12
584,12
585,12
586,12
587,12
588,12
589,12
590,12
591,12
592,12
593,12
594,12
595,12
596,12
597,12
598,12
599,12
600,12
601,12
602,12
603,12
604,12
605,12
606,12
607,12
608,12
609,12
610,12
611,12
612,12
613,12
614,12
615,12
616,12
617,12
618,12
619,12
620,12
621,12
622,12
623,12
624,13
625,13
626,13
627,13
628,13
629,13
630,13
631,13
632,13
633,13
634,13
635,13
636,13
637,13
638,13
639,13
640,13
641,13
642,13
643,13
644,13
645,13
646,13
647,13
648,13
649,13
650,13
651,13
652,13
653,13
654,13
655,13
656,13
657,13
658,13
659,13
660,13
661,13
662,13
663,13
664,13
665,13
666,13
667,13
668,13
669,13
670,13
671,13
672,14
673,14
674,14
675,14
676,14
677,14
678,14
679,14
680,14
681,14
682,14
683,14
684,14
685,14
686,14
687,14
688,14
689,14
690,14
691,14
692,14
693,14
694,14
695,14
696,14
697,14
698,14
699,14
700,14
701,14
702,14
703,14
704,14
705,14
706,14
707,14
708,14
709,14
710,14
711,14
712,14
713,14
714,14
715,14
716,14
717,14
718,14
719,14
720,15
721,15
722,15
723,15
724,15
725,15
726,15
727,15
728,15
729,15
730,15
731,15
732,15
733,15
734,15
735,15
736,15
737,15
738,15
739,15
740,15
741,15
742,15
743,15
744,15
745,15
746,15
747,15
748,15
749,15
750,15
751,15
752,15
753,15
754,15
755,15
756,15
757,15
758,15
759,15
760,15
761,15
762,15
763,15
764,15
765,15
766,15
767,15
768,16
769,16
770,16
771,16
772,16
773,16
774,16
775,16
776,16
777,16
778,16
779,16
780,16
781,16
782,16
783,16
784,16
785,16
786,16
787,16
788,16
789,16
790,16
791,16
792,16
793,16
794,16
795,16
796,16
797,16
798,16
799,16
800,16
801,16
802,16
803,16
804,16
805,16
806,16
807,16
808,16
809,16
810,16
811,16
812,16
813,16
814,16
815,16
816,17
817,17
818,17
819,17
820,17
821,17
822,17
823,17
824,17
825,17
826,17
827,17
828,17
829,17
830,17
831,17
832,17
833,17
834,17
835,17
836,17
837,17
838,17
839,17
840,17
841,17
842,17
843,17
844,17
845,17
846,17
847,17
848,17
849,17
850,17
851,17
852,17
853,17
854,17
855,17
856,17
857,17
858,17
859,17
860,17
861,17
862,17
863,17
864,18
865,18
866,18
867,18
868,18
869,18
870,18
871,18
872,18
873,18
874,18
875,18
876,18
877,18
878,18
879,18
880,18
881,18
882,18
883,18
884,18
885,18
886,18
887,18
888,18
889,18
890,18
891,18
892,18
893,18
894,18
895,18
896,18
897,18
898,18
899,18
900,18
901,18
902,18
903,18
904,18
905,18
906,18
907,18
908,18
909,18
910,18
911,18
912,19
913,19
914,19
915,19
916,19
917,19
918,19
919,19
920,19
921,19
922,19
923,19
924,19
925,19
926,19
927,19
928,19
929,19
930,19
931,19
932,19
933,19
934,19
935,19
936,19
937,19
938,19
939,19
940,19
941,19
942,19
943,19
944,19
945,19
946,19
947,19
948,19
949,19
950,19
951,19
952,19
953,19
954,19
955,19
956,19
957,19
958,19
959,19
960,20
961,20
962,20
963,20
964,20
965,20
966,20
967,20
968,20
969,20
970,20
971,20
972,20
973,20
974,20
975,20
976,20
977,20
978,20
979,20
980,20
981,20
982,20
983,20
984,20
985,20
986,20
987,20
988,20
989,20
990,20
991,20
992,20
993,20
994,20
995,20
996,20
997,20
998,20
999,20
1000,20
1001,20
1002,20
1003,20
1004,20
1005,20
1006,20
1007,20
1008,21
1009,21
1010,21
1011,21
1012,21
1013,21
1014,21
1015,21
1016,21
1017,21
1018,21
1019,21
1020,21
1021,21
1022,21
1023,21
1024,21
1025,21
1026,21
1027,21
1028,21
1029,21
1030,21
1031,21
1032,21
1033,21
1034,21
1035,21
1036,21
1037,21
1038,21
1039,21
1040,21
1041,21
1042,21
1043,21
1044,21
1045,21
1046,21
1047,21
1048,21
1049,21
1050,21
1051,21
1052,21
1053,21
1054,21
1055,21
1056,22
1057,22
1058,22
1059,22
1060,22
1061,22
1062,22
1063,22
1064,22
1065,22
1066,22
1067,22
1068,22
1069,22
1070,22
1071,22
1072,22
1073,22
1074,22
1075,22
1076,22
1077,22
1078,22
1079,22
1080,22
1081,22
1082,22
1083,22
1084,22
1085,22
1086,22
1087,22
1088,22
1089,22
1090,22
1091,22
1092,22
1093,22
1094,22
1095,22
1096,22
1097,22
1098,22
1099,22
1100,22
1101,22
1102,22
1103,22
1104,23
1105,23
1106,23
1107,23
1108,23
1109,23
1110,23
1111,23
1112,23
1113,23
1114,23
1115,23
1116,23
1117,23
1118,23
1119,23
1120,23
1121,23
1122,23
1123,23
1124,23
1125,23
1126,23
1127,23
1128,23
1129,23
1130,23
1131,23
1132,23
1133,23
1134,23
1135,23
1136,23
1137,23
1138,23
1139,23
1140,23
1141,23
1142,23
1143,23
1144,23
1145,23
1146,23
1147,23
1148,23
1149,23
1150,23
1151,23
1152,24
1153,24
1154,24
1155,24
1156,24
1157,24
1158,24
1159,24
1160,24
1161,24
1162,24
1163,24
1164,24
1165,24
1166,24
1167,24
1168,24
1169,24
1170,24
1171,24
1172,24
1173,24
1174,24
1175,24
1176,24
1177,24
1178,24
1179,24
1180,24
1181,24
1182,24
1183,24
1184,24
1185,24
1186,24
1187,24
1188,24
1189,24
1190,24
1191,24
1192,24
1193,24
1194,24
1195,24
1196,24
1197,24
1198,24
1199,24
1200,25
1201,25
1202,25
1203,25
1204,25
1205,25
1206,25
1207,25
1208,25
1209,25
1210,25
1211,25
1212,25
1213,25
1214,25
1215,25
1216,25
1217,25
1218,25
1219,25
1220,25
1221,25
1222,25
1223,25
1224,25
1225,25
1226,25
1227,25
1228,25
1229,25
1230,25
1231,25
1232,25
1233,25
1234,25
1235,25
1236,25
1237,25
1238,25
1239,25
1240,25
1241,25
1242,25
1243,25
1244,25
1245,25
1246,25
1247,25
1248,26
1249,26
1250,26
1251,26
1252,26
1253,26
1254,26
1255,26
1256,26
1257,26
1258,26
1259,26
1260,26
1261,26
1262,26
1263,26
1264,26
1265,26
1266,26
1267,26
1268,26
1269,26
1270,26
1271,26
1272,26
1273,26
1274,26
1275,26
1276,26
1277,26
1278,26
1279,26
1280,26
1281,26
1282,26
1283,26
1284,26
1285,26
1286,26
1287,26
1288,26
1289,26
1290,26
1291,26
1292,26
1293,26
1294,26
1295,26
1296,27
1297,27
1298,27
1299,27
1300,27
1301,27
1302,27
1303,27
1304,27
1305,27
1306,27
1307,27
1308,27
1309,27
1310,27
1311,27
1312,27
1313,27
1314,27
1315,27
1316,27
1317,27
1318,27
1319,27
1320,27
1321,27
1322,27
1323,27
1324,27
1325,27
1326,27
1327,27
1328,27
1329,27
1330,27
1331,27
1332,27
1333,27
1334,27
1335,27
1336,27
1337,27
1338,27
1339,27
1340,27
1341,27
1342,27
1343,27
1344,28
1345,28
1346,28
1347,28
1348,28
1349,28
1350,28
1351,28
1352,28
1353,28
1354,28
1355,28
1356,28
1357,28
1358,28
1359,28
1360,28
1361,28
1362,28
1363,28
1364,28
1365,28
1366,28
1367,28
1368,28
1369,28
1370,28
1371,28
1372,28
1373,28
1374,28
1375,28
1376,28
1377,28
1378,28
1379,28
1380,28
1381,28
1382,28
1383,28
1384,28
1385,28
1386,28
1387,28
1388,28
1389,28
1390,28
1391,28
1392,29
1393,29
1394,29
1395,29
1396,29
1397,29
1398,29
1399,29
1400,29
1401,29
1402,29
1403,29
1404,29
1405,29
1406,29
1407,29
1408,29
1409,29
1410,29
1411,29
1412,29
1413,29
1414,29
1415,29
1416,29
1417,29
1418,29
1419,29
1420,29
1421,29
1422,29
1423,29
1424,29
1425,29
1426,29
1427,29
1428,29
1429,29
1430,29
1431,29
1432,29
1433,29
1434,29
1435,29
1436,29
1437,29
1438,29
1439,29
1440,30
1441,30
1442,30
1443,30
1444,30
1445,30
1446,30
1447,30
1448,30
1449,30
1450,30
1451,30
1452,30
1453,30
1454,30
1455,30
1456,30
1457,30
1458,30
1459,30
1460,30
1461,30
1462,30
1463,30
1464,30
1465,30
1466,30
1467,30
1468,30
1469,30
1470,30
1471,30
1472,30
1473,30
1474,30
1475,30
1476,30
1477,30
1478,30
1479,30
1480,30
1481,30
1482,30
1483,30
1484,30
1485,30
1486,30
1487,30
1488,31
1489,31
1490,31
1491,31
1492,31
1493,31
1494,31
1495,31
1496,31
1497,31
1498,31
1499,31
1500,31
1501,31
1502,31
1503,31
1504,31
1505,31
1506,31
1507,31
1508,31
1509,31
1510,31
1511,31
1512,31
1513,31
1514,31
1515,31
1516,31
1517,31
1518,31
1519,31
1520,31
1521,31
1522,31
1523,31
1524,31
1525,31
1526,31
1527,31
1528,31
1529,31
1530,31
1531,31
1532,31
1533,31
1534,31
1535,31
1536,32
1537,32
1538,32
1539,32
1540,32
1541,32
1542,32
1543,32
1544,32
1545,32
1546,32
1547,32
1548,32
1549,32
1550,32
1551,32
1552,32
1553,32
1554,32
1555,32
1556,32
1557,32
1558,32
1559,32
1560,32
1561,32
1562,32
1563,32
1564,32
1565,32
1566,32
1567,32
1568,32
1569,32
1570,32
1571,32
1572,32
1573,32
1574,32
1575,32
1576,32
1577,32
1578,32
1579,32
1580,32
1581,32
1582,32
1583,32
1584,33
1585,33
1586,33
1587,33
1588,33
1589,33
1590,33
1591,33
1592,33
1593,33
1594,33
1595,33
1596,33
1597,33
1598,33
1599,33
1600,33
1601,33
1602,33
1603,33
1604,33
1605,33
1606,33
1607,33
1608,33
1609,33
1610,33
1611,33
1612,33
1613,33
1614,33
1615,33
1616,33
1617,33
1618,33
1619,33
1620,33
1621,33
1622,33
1623,33
1624,33
1625,33
1626,33
1627,33
1628,33
1629,33
1630,33
1631,33
1632,34
1633,34
1634,34
1635,34
1636,34
1637,34
1638,34
1639,34
1640,34
1641,34
1642,34
1643,34
1644,34
1645,34
1646,34
1647,34
1648,34
1649,34
1650,34
1651,34
1652,34
1653,34
1654,34
1655,34
1656,34
1657,34
1658,34
1659,34
1660,34
1661,34
1662,34
1663,34
1664,34
1665,34
1666,34
1667,34
1668,34
1669,34
1670,34
1671,34
1672,34
1673,34
1674,34
1675,34
1676,34
1677,34
1678,34
1679,34
1680,35
1681,35
1682,35
1683,35
1684,35
1685,35
1686,35
1687,35
1688,35
1689,35
1690,35
1691,35
1692,35
1693,35
1694,35
1695,35
1696,35
1697,35
1698,35
1699,35
1700,35
1701,35
1702,35
1703,35
1704,35
1705,35
1706,35
1707,35
1708,35
1709,35
1710,35
1711,35
1712,35
1713,35
1714,35
1715,35
1716,35
1717,35
1718,35
1719,35
1720,35
1721,35
1722,35
1723,35
1724,35
1725,35
1726,35
1727,35
1728,36
1729,36
1730,36
1731,36
1732,36
1733,36
1734,36
1735,36
1736,36
1737,36
1738,36
1739,36
1740,36
1741,36
1742,36
1743,36
1744,36
1745,36
1746,36
1747,36
1748,36
1749,36
1750,36
1751,36
1752,36
1753,36
1754,36
1755,36
1756,36
1757,36
1758,36
1759,36
1760,36
1761,36
1762,36
1763,36
1764,36
1765,36
1766,36
1767,36
1768,36
1769,36
1770,36
1771,36
1772,36
1773,36
1774,36
1775,36
1776,37
1777,37
1778,37
1779,37
1780,37
1781,37
1782,37
1783,37
1784,37
1785,37
1786,37
1787,37
1788,37
1789,37
1790,37
1791,37
1792,37
1793,37
1794,37
1795,37
1796,37
1797,37
1798,37
1799,37
1800,37
1801,37
1802,37
1803,37
1804,37
1805,37
1806,37
1807,37
1808,37
1809,37
1810,37
1811,37
1812,37
1813,37
1814,37
1815,37
1816,37
1817,37
1818,37
1819,37
1820,37
1821,37
1822,37
1823,37
1824,38
1825,38
1826,38
1827,38
1828,38
1829,38
1830,38
1831,38
1832,38
1833,38
1834,38
1835,38
1836,38
1837,38
1838,38
1839,38
1840,38
1841,38
1842,38
1843,38
1844,38
1845,38
1846,38
1847,38
1848,38
1849,38
1850,38
1851,38
1852,38
1853,38
1854,38
1855,38
1856,38
1857,38
1858,38
1859,38
1860,38
1861,38
1862,38
1863,38
1864,38
1865,38
1866,38
1867,38
1868,38
1869,38
1870,38
1871,38
1872,39
1873,39
1874,39
1875,39
1876,39
1877,39
1878,39
1879,39
1880,39
1881,39
1882,39
1883,39
1884,39
1885,39
1886,39
1887,39
1888,39
1889,39
1890,39
1891,39
1892,39
1893,39
1894,39
1895,39
1896,39
1897,39
1898,39
1899,39
1900,39
1901,39
1902,39
1903,39
1904,39
1905,39
1906,39
1907,39
1908,39
1909,39
1910,39
1911,39
1912,39
1913,39
1914,39
1915,39
1916,39
1917,39
1918,39
1919,39
1920,40
1921,40
1922,40
1923,40
1924,40
1925,40
1926,40
1927,40
1928,40
1929,40
1930,40
1931,40
1932,40
1933,40
1934,40
1935,40
1936,40
1937,40
1938,40
1939,40
1940,40
1941,40
1942,40
1943,40
1944,40
1945,40
1946,40
1947,40
1948,40
1949,40
1950,40
1951,40
1952,40
1953,40
1954,40
1955,40
1956,40
1957,40
1958,40
1959,40
1960,40
1961,40
1962,40
1963,40
1964,40
1965,40
1966,40
1967,40
1968,41
1969,41
1970,41
1971,41
1972,41
1973,41
1974,41
1975,41
1976,41
1977,41
1978,41
1979,41
1980,41
1981,41
1982,41
1983,41
1984,41
1985,41
1986,41
1987,41
1988,41
1989,41
1990,41
1991,41
1992,41
1993,41
1994,41
1995,41
1996,41
1997,41
1998,41
1999,41
2000,41
2001,41
2002,41
2003,41
2004,41
2005,41
2006,41
2007,41
2008,41
2009,41
2010,41
2011,41
2012,41
2013,41
2014,41
2015,41
2016,42
2017,42
2018,42
2019,42
2020,42
2021,42
2022,42
2023,42
2024,42
2025,42
2026,42
2027,42
2028,42
2029,42
2030,42
2031,42
2032,42
2033,42
2034,42
2035,42
2036,42
2037,42
2038,42
2039,42
2040,42
2041,42
2042,42
2043,42
2044,42
2045,42
2046,42
2047,42
2048,42
2049,42
2050,42
2051,42
2052,42
2053,42
2054,42
2055,42
2056,42
2057,42
2058,42
2059,42
2060,42
2061,42
2062,42
2063,42
2064,43
2065,43
2066,43
2067,43
2068,43
2069,43
2070,43
2071,43
2072,43
2073,43
2074,43
2075,43
2076,43
2077,43
2078,43
2079,43
2080,43
2081,43
2082,43
2083,43
2084,43
2085,43
2086,43
2087,43
2088,43
2089,43
2090,43
2091,43
2092,43
2093,43
2094,43
2095,43
2096,43
2097,43
2098,43
2099,43
2100,43
2101,43
2102,43
2103,43
2104,43
2105,43
2106,43
2107,43
2108,43
2109,43
2110,43
2111,43
2112,44
2113,44
2114,44
2115,44
2116,44
2117,44
2118,44
2119,44
2120,44
2121,44
2122,44
2123,44
2124,44
2125,44
2126,44
2127,44
2128,44
2129,44
2130,44
2131,44
2132,44
2133,44
2134,44
2135,44
2136,44
2137,44
2138,44
2139,44
2140,44
2141,44
2142,44
2143,44
2144,44
2145,44
2146,44
2147,44
2148,44
2149,44
2150,44
2151,44
2152,44
2153,44
2154,44
2155,44
2156,44
2157,44
2158,44
2159,44
2160,45
2161,45
2162,45
2163,45
2164,45
2165,45
2166,45
2167,45
2168,45
2169,45
2170,45
2171,45
2172,45
2173,45
2174,45
2175,45
2176,45
2177,45
2178,45
2179,45
2180,45
2181,45
2182,45
2183,45
2184,45
2185,45
2186,45
2187,45
2188,45
2189,45
2190,45
2191,45
2192,45
2193,45
2194,45
2195,45
2196,45
2197,45
2198,45
2199,45
2200,45
2201,45
2202,45
2203,45
2204,45
2205,45
2206,45
2207,45
2208,46
2209,46
2210,46
2211,46
2212,46
2213,46
2214,46
2215,46
2216,46
2217,46
2218,46
2219,46
2220,46
2221,46
2222,46
2223,46
2224,46
2225,46
2226,46
2227,46
2228,46
2229,46
2230,46
2231,46
2232,46
2233,46
2234,46
2235,46
2236,46
2237,46
2238,46
2239,46
2240,46
2241,46
2242,46
2243,46
2244,46
2245,46
2246,46
2247,46
2248,46
2249,46
2250,46
2251,46
2252,46
2253,46
2254,46
2255,46
2256,47
2257,47
2258,47
2259,47
2260,47
2261,47
2262,47
2263,47
2264,47
2265,47
2266,47
2267,47
2268,47
2269,47
2270,47
2271,47
2272,47
2273,47
2274,47
2275,47
2276,47
2277,47
2278,47
2279,47
2280,47
2281,47
2282,47
2283,47
2284,47
2285,47
2286,47
2287,47
2288,47
2289,47
2290,47
2291,47
2292,47
2293,47
2294,47
2295,47
2296,47
2297,47
2298,47
2299,47
2300,47
2301,47
2302,47
2303,47
2304,48
2305,48
2306,48
2307,48
2308,48
2309,48
2310,48
2311,48
2312,48
2313,48
2314,48
2315,48
2316,48
2317,48
2318,48
2319,48
2320,48
2321,48
2322,48
2323,48
2324,48
2325,48
2326,48
2327,48
2328,48
2329,48
2330,48
2331,48
2332,48
2333,48
2334,48
2335,48
2336,48
2337,48
2338,48
2339,48
2340,48
2341,48
2342,48
2343,48
2344,48
2345,48
2346,48
2347,48
2348,48
2349,48
2350,48
2351,48
2352,49
2353,49
2354,49
2355,49
2356,49
2357,49
2358,49
2359,49
2360,49
2361,49
2362,49
2363,49
2364,49
2365,49
2366,49
2367,49
2368,49
2369,49
2370,49
2371,49
2372,49
2373,49
2374,49
2375,49
2376,49
2377,49
2378,49
2379,49
2380,49
2381,49
2382,49
2383,49
2384,49
2385,49
2386,49
2387,49
2388,49
2389,49
2390,49
2391,49
2392,49
2393,49
2394,49
2395,49
2396,49
2397,49
2398,49
2399,49
2400,50
2401,50
2402,50
2403,50
2404,50
2405,50
2406,50
2407,50
2408,50
2409,50
2410,50
2411,50
2412,50
2413,50
2414,50
2415,50
2416,50
2417,50
2418,50
2419,50
2420,50
2421,50
2422,50
2423,50
2424,50
2425,50
2426,50
2427,50
2428,50
2429,50
2430,50
2431,50
2432,50
2433,50
2434,50
2435,50
2436,50
2437,50
2438,50
2439,50
2440,50
2441,50
2442,50
2443,50
2444,50
2445,50
2446,50
2447,50
2448,51
2449,51
2450,51
2451,51
2452,51
2453,51
2454,51
2455,51
2456,51
2457,51
2458,51
2459,51
2460,51
2461,51
2462,51
2463,51
2464,51
2465,51
2466,51
2467,51
2468,51
2469,51
2470,51
2471,51
2472,51
2473,51
2474,51
2475,51
2476,51
2477,51
2478,51
2479,51
2480,51
2481,51
2482,51
2483,51
2484,51
2485,51
2486,51
2487,51
2488,51
2489,51
2490,51
2491,51
2492,51
2493,51
2494,51
2495,51
2496,52
2497,52
2498,52
2499,52
2500,52
2501,52
2502,52
2503,52
2504,52
2505,52
2506,52
2507,52
2508,52
2509,52
2510,52
2511,52
2512,52
2513,52
2514,52
2515,52
2516,52
2517,52
2518,52
2519,52
2520,52
2521,52
2522,52
2523,52
2524,52
2525,52
2526,52
2527,52
2528,52
2529,52
2530,52
2531,52
2532,52
2533,52
2534,52
2535,52
2536,52
2537,52
2538,52
2539,52
2540,52
2541,52
2542,52
2543,52
2544,53
2545,53
2546,53
2547,53
2548,53
2549,53
2550,53
2551,53
2552,53
2553,53
2554,53
2555,53
2556,53
2557,53
2558,53
2559,53
2560,53
2561,53
2562,53
2563,53
2564,53
2565,53
2566,53
2567,53
2568,53
2569,53
2570,53
2571,53
2572,53
2573,53
2574,53
2575,53
2576,53
2577,53
2578,53
2579,53
2580,53
2581,53
2582,53
2583,53
2584,53
2585,53
2586,53
2587,53
2588,53
2589,53
2590,53
2591,53
2592,54
2593,54
2594,54
2595,54
2596,54
2597,54
2598,54
2599,54
2600,54
2601,54
2602,54
2603,54
2604,54
2605,54
2606,54
2607,54
2608,54
2609,54
2610,54
2611,54
2612,54
2613,54
2614,54
2615,54
2616,54
2617,54
2618,54
2619,54
2620,54
2621,54
2622,54
2623,54
2624,54
2625,54
2626,54
2627,54
2628,54
2629,54
2630,54
2631,54
2632,54
2633,54
2634,54
2635,54
2636,54
2637,54
2638,54
2639,54
2640,55
2641,55
2642,55
2643,55
2644,55
2645,55
2646,55
2647,55
2648,55
2649,55
2650,55
2651,55
2652,55
2653,55
2654,55
2655,55
2656,55
2657,55
2658,55
2659,55
2660,55
2661,55
2662,55
2663,55
2664,55
2665,55
2666,55
2667,55
2668,55
2669,55
2670,55
2671,55
2672,55
2673,55
2674,55
2675,55
2676,55
2677,55
2678,55
2679,55
2680,55
2681,55
2682,55
2683,55
2684,55
2685,55
2686,55
2687,55
2688,56
2689,56
2690,56
2691,56
2692,56
2693,56
2694,56
2695,56
2696,56
2697,56
2698,56
2699,56
2700,56
2701,56
2702,56
2703,56
2704,56
2705,56
2706,56
2707,56
2708,56
2709,56
2710,56
2711,56
2712,56
2713,56
2714,56
2715,56
2716,56
2717,56
2718,56
2719,56
2720,56
2721,56
2722,56
2723,56
2724,56
2725,56
2726,56
2727,56
2728,56
2729,56
2730,56
2731,56
2732,56
2733,56
2734,56
2735,56
2736,57
2737,57
2738,57
2739,57
2740,57
2741,57
2742,57
2743,57
2744,57
2745,57
2746,57
2747,57
2748,57
2749,57
2750,57
2751,57
2752,57
2753,57
2754,57
2755,57
2756,57
2757,57
2758,57
2759,57
2760,57
2761,57
2762,57
2763,57
2764,57
2765,57
2766,57
2767,57
2768,57
2769,57
2770,57
2771,57
2772,57
2773,57
2774,57
2775,57
2776,57
2777,57
2778,57
2779,57
2780,57
2781,57
2782,57
2783,57
2784,58
2785,58
2786,58
2787,58
2788,58
2789,58
2790,58
2791,58
2792,58
2793,58
2794,58
2795,58
2796,58
2797,58
2798,58
2799,58
2800,58
2801,58
2802,58
2803,58
2804,58
2805,58
2806,58
2807,58
2808,58
2809,58
2810,58
2811,58
2812,58
2813,58
2814,58
2815,58
2816,58
2817,58
2818,58
2819,58
2820,58
2821,58
2822,58
2823,58
2824,58
2825,58
2826,58
2827,58
2828,58
2829,58
2830,58
2831,58
2832,59
2833,59
2834,59
2835,59
2836,59
2837,59
2838,59
2839,59
2840,59
2841,59
2842,59
2843,59
2844,59
2845,59
2846,59
2847,59
2848,59
2849,59
2850,59
2851,59
2852,59
2853,59
2854,59
2855,59
2856,59
2857,59
2858,59
2859,59
2860,59
2861,59
2862,59
2863,59
2864,59
2865,59
2866,59
2867,59
2868,59
2869,59
2870,59
2871,59
2872,59
2873,59
2874,59
2875,59
2876,59
2877,59
2878,59
2879,59
2880,60
2881,60
2882,60
2883,60
2884,60
2885,60
2886,60
2887,60
2888,60
2889,60
2890,60
2891,60
2892,60
2893,60
2894,60
2895,60
2896,60
2897,60
2898,60
2899,60
2900,60
2901,60
2902,60
2903,60
2904,60
2905,60
2906,60
2907,60
2908,60
2909,60
2910,60
2911,60
2912,60
2913,60
2914,60
2915,60
2916,60
2917,60
2918,60
2919,60
2920,60
2921,60
2922,60
2923,60
2924,60
2925,60
2926,60
2927,60
2928,61
2929,61
2930,61
2931,61
2932,61
2933,61
2934,61
2935,61
2936,61
2937,61
2938,61
2939,61
2940,61
2941,61
2942,61
2943,61
2944,61
2945,61
2946,61
2947,61
2948,61
2949,61
2950,61
2951,61
2952,61
2953,61
2954,61
2955,61
2956,61
2957,61
2958,61
2959,61
2960,61
2961,61
2962,61
2963,61
2964,61
2965,61
2966,61
2967,61
2968,61
2969,61
2970,61
2971,61
2972,61
2973,61
2974,61
2975,61
2976,62
2977,62
2978,62
2979,62
2980,62
2981,62
2982,62
2983,62
2984,62
2985,62
2986,62
2987,62
2988,62
2989,62
2990,62
2991,62
2992,62
2993,62
2994,62
2995,62
2996,62
2997,62
2998,62
2999,62
3000,62
3001,62
3002,62
3003,62
3004,62
3005,62
3006,62
3007,62
3008,62
3009,62
3010,62
3011,62
3012,62
3013,62
3014,62
3015,62
3016,62
3017,62
3018,62
3019,62
3020,62
3021,62
3022,62
3023,62
3024,63
3025,63
3026,63
3027,63
3028,63
3029,63
3030,63
3031,63
3032,63
3033,63
3034,63
3035,63
3036,63
3037,63
3038,63
3039,63
3040,63
3041,63
3042,63
3043,63
3044,63
3045,63
3046,63
3047,63
3048,63
3049,63
3050,63
3051,63
3052,63
3053,63
3054,63
3055,63
3056,63
3057,63
3058,63
3059,63
3060,63
3061,63
3062,63
3063,63
3064,63
3065,63
3066,63
3067,63
3068,63
3069,63
3070,63
3071,63
3072,64
3073,64
3074,64
3075,64
3076,64
3077,64
3078,64
3079,64
3080,64
3081,64
3082,64
3083,64
3084,64
3085,64
3086,64
3087,64
3088,64
3089,64
3090,64
3091,64
3092,64
3093,64
3094,64
3095,64
3096,64
3097,64
3098,64
3099,64
3100,64
3101,64
3102,64
3103,64
3104,64
3105,64
3106,64
3107,64
3108,64
3109,64
3110,64
3111,64
3112,64
3113,64
3114,64
3115,64
3116,64
3117,64
3118,64
3119,64
3120,65
3121,65
3122,65
3123,65
3124,65
3125,65
3126,65
3127,65
3128,65
3129,65
3130,65
3131,65
3132,65
3133,65
3134,65
3135,65
3136,65
3137,65
3138,65
3139,65
3140,65
3141,65
3142,65
3143,65
3144,65
3145,65
3146,65
3147,65
3148,65
3149,65
3150,65
3151,65
3152,65
3153,65
3154,65
3155,65
3156,65
3157,65
3158,65
3159,65
3160,65
3161,65
3162,65
3163,65
3164,65
3165,65
3166,65
3167,65
3168,66
3169,66
3170,66
3171,66
3172,66
3173,66
3174,66
3175,66
3176,66
3177,66
3178,66
3179,66
3180,66
3181,66
3182,66
3183,66
3184,66
3185,66
3186,66
3187,66
3188,66
3189,66
3190,66
3191,66
3192,66
3193,66
3194,66
3195,66
3196,66
3197,66
3198,66
3199,66
3200,66
3201,66
3202,66
3203,66
3204,66
3205,66
3206,66
3207,66
3208,66
3209,66
3210,66
3211,66
3212,66
3213,66
3214,66
3215,66
3216,67
3217,67
3218,67
3219,67
3220,67
3221,67
3222,67
3223,67
3224,67
3225,67
3226,67
3227,67
3228,67
3229,67
3230,67
3231,67
3232,67
3233,67
3234,67
3235,67
3236,67
3237,67
3238,67
3239,67
3240,67
3241,67
3242,67
3243,67
3244,67
3245,67
3246,67
3247,67
3248,67
3249,67
3250,67
3251,67
3252,67
3253,67
3254,67
3255,67
3256,67
3257,67
3258,67
3259,67
3260,67
3261,67
3262,67
3263,67
3264,68
3265,68
3266,68
3267,68
3268,68
3269,68
3270,68
3271,68
3272,68
3273,68
3274,68
3275,68
3276,68
3277,68
3278,68
3279,68
3280,68
3281,68
3282,68
3283,68
3284,68
3285,68
3286,68
3287,68
3288,68
3289,68
3290,68
3291,68
3292,68
3293,68
3294,68
3295,68
3296,68
3297,68
3298,68
3299,68
3300,68
3301,68
3302,68
3303,68
3304,68
3305,68
3306,68
3307,68
3308,68
3309,68
3310,68
3311,68
3312,69
3313,69
3314,69
3315,69
3316,69
3317,69
3318,69
3319,69
3320,69
3321,69
3322,69
3323,69
3324,69
3325,69
3326,69
3327,69
3328,69
3329,69
3330,69
3331,69
3332,69
3333,69
3334,69
3335,69
3336,69
3337,69
3338,69
3339,69
3340,69
3341,69
3342,69
3343,69
3344,69
3345,69
3346,69
3347,69
3348,69
3349,69
3350,69
3351,69
3352,69
3353,69
3354,69
3355,69
3356,69
3357,69
3358,69
3359,69
3360,70
3361,70
3362,70
3363,70
3364,70
3365,70
3366,70
3367,70
3368,70
3369,70
3370,70
3371,70
3372,70
3373,70
3374,70
3375,70
3376,70
3377,70
3378,70
3379,70
3380,70
3381,70
3382,70
3383,70
3384,70
3385,70
3386,70
3387,70
3388,70
3389,70
3390,70
3391,70
3392,70
3393,70
3394,70
3395,70
3396,70
3397,70
3398,70
3399,70
3400,70
3401,70
3402,70
3403,70
3404,70
3405,70
3406,70
3407,70
3408,71
3409,71
3410,71
3411,71
3412,71
3413,71
3414,71
3415,71
3416,71
3417,71
3418,71
3419,71
3420,71
3421,71
3422,71
3423,71
3424,71
3425,71
3426,71
3427,71
3428,71
3429,71
3430,71
3431,71
3432,71
3433,71
3434,71
3435,71
3436,71
3437,71
3438,71
3439,71
3440,71
3441,71
3442,71
3443,71
3444,71
3445,71
3446,71
3447,71
3448,71
3449,71
3450,71
3451,71
3452,71
3453,71
3454,71
3455,71
3456,72
3457,72
3458,72
3459,72
3460,72
3461,72
3462,72
3463,72
3464,72
3465,72
3466,72
3467,72
3468,72
3469,72
3470,72
3471,72
3472,72
3473,72
3474,72
3475,72
3476,72
3477,72
3478,72
3479,72
3480,72
3481,72
3482,72
3483,72
3484,72
3485,72
3486,72
3487,72
3488,72
3489,72
3490,72
3491,72
3492,72
3493,72
3494,72
3495,72
3496,72
3497,72
3498,72
3499,72
3500,72
3501,72
3502,72
3503,72
3504,73
3505,73
3506,73
3507,73
3508,73
3509,73
3510,73
3511,73
3512,73
3513,73
3514,73
3515,73
3516,73
3517,73
3518,73
3519,73
3520,73
3521,73
3522,73
3523,73
3524,73
3525,73
3526,73
3527,73
3528,73
3529,73
3530,73
3531,73
3532,73
3533,73
3534,73
3535,73
3536,73
3537,73
3538,73
3539,73
3540,73
3541,73
3542,73
3543,73
3544,73
3545,73
3546,73
3547,73
3548,73
3549,73
3550,73
3551,73
3552,74
3553,74
3554,74
3555,74
3556,74
3557,74
3558,74
3559,74
3560,74
3561,74
3562,74
3563,74
3564,74
3565,74
3566,74
3567,74
3568,74
3569,74
3570,74
3571,74
3572,74
3573,74
3574,74
3575,74
3576,74
3577,74
3578,74
3579,74
3580,74
3581,74
3582,74
3583,74
3584,74
3585,74
3586,74
3587,74
3588,74
3589,74
3590,74
3591,74
3592,74
3593,74
3594,74
3595,74
3596,74
3597,74
3598,74
3599,74
3600,75
3601,75
3602,75
3603,75
3604,75
3605,75
3606,75
3607,75
3608,75
3609,75
3610,75
3611,75
3612,75
3613,75
3614,75
3615,75
3616,75
3617,75
3618,75
3619,75
3620,75
3621,75
3622,75
3623,75
3624,75
3625,75
3626,75
3627,75
3628,75
3629,75
3630,75
3631,75
3632,75
3633,75
3634,75
3635,75
3636,75
3637,75
3638,75
3639,75
3640,75
3641,75
3642,75
3643,75
3644,75
3645,75
3646,75
3647,75
3648,76
3649,76
3650,76
3651,76
3652,76
3653,76
3654,76
3655,76
3656,76
3657,76
3658,76
3659,76
3660,76
3661,76
3662,76
3663,76
3664,76
3665,76
3666,76
3667,76
3668,76
3669,76
3670,76
3671,76
3672,76
3673,76
3674,76
3675,76
3676,76
3677,76
3678,76
3679,76
3680,76
3681,76
3682,76
3683,76
3684,76
3685,76
3686,76
3687,76
3688,76
3689,76
3690,76
3691,76
3692,76
3693,76
3694,76
3695,76
3696,77
3697,77
3698,77
3699,77
3700,77
3701,77
3702,77
3703,77
3704,77
3705,77
3706,77
3707,77
3708,77
3709,77
3710,77
3711,77
3712,77
3713,77
3714,77
3715,77
3716,77
3717,77
3718,77
3719,77
3720,77
3721,77
3722,77
3723,77
3724,77
3725,77
3726,77
3727,77
3728,77
3729,77
3730,77
3731,77
3732,77
3733,77
3734,77
3735,77
3736,77
3737,77
3738,77
3739,77
3740,77
3741,77
3742,77
3743,77
3744,78
3745,78
3746,78
3747,78
3748,78
3749,78
3750,78
3751,78
3752,78
3753,78
3754,78
3755,78
3756,78
3757,78
3758,78
3759,78
3760,78
3761,78
3762,78
3763,78
3764,78
3765,78
3766,78
3767,78
3768,78
3769,78
3770,78
3771,78
3772,78
3773,78
3774,78
3775,78
3776,78
3777,78
3778,78
3779,78
3780,78
3781,78
3782,78
3783,78
3784,78
3785,78
3786,78
3787,78
3788,78
3789,78
3790,78
3791,78
3792,79
3793,79
3794,79
3795,79
3796,79
3797,79
3798,79
3799,79
3800,79
3801,79
3802,79
3803,79
3804,79
3805,79
3806,79
3807,79
3808,79
3809,79
3810,79
3811,79
3812,79
3813,79
3814,79
3815,79
3816,79
3817,79
3818,79
3819,79
3820,79
3821,79
3822,79
3823,79
3824,79
3825,79
3826,79
3827,79
3828,79
3829,79
3830,79
3831,79
3832,79
3833,79
3834,79
3835,79
3836,79
3837,79
3838,79
3839,79
3840,80
3841,80
3842,80
3843,80
3844,80
3845,80
3846,80
3847,80
3848,80
3849,80
3850,80
3851,80
3852,80
3853,80
3854,80
3855,80
3856,80
3857,80
3858,80
3859,80
3860,80
3861,80
3862,80
3863,80
3864,80
3865,80
3866,80
3867,80
3868,80
3869,80
3870,80
3871,80
3872,80
3873,80
3874,80
3875,80
3876,80
3877,80
3878,80
3879,80
3880,80
3881,80
3882,80
3883,80
3884,80
3885,80
3886,80
3887,80
3888,81
3889,81
3890,81
3891,81
3892,81
3893,81
3894,81
3895,81
3896,81
3897,81
3898,81
3899,81
3900,81
3901,81
3902,81
3903,81
3904,81
3905,81
3906,81
3907,81
3908,81
3909,81
3910,81
3911,81
3912,81
3913,81
3914,81
3915,81
3916,81
3917,81
3918,81
3919,81
3920,81
3921,81
3922,81
3923,81
3924,81
3925,81
3926,81
3927,81
3928,81
3929,81
3930,81
3931,81
3932,81
3933,81
3934,81
3935,81
3936,82
3937,82
3938,82
3939,82
3940,82
3941,82
3942,82
3943,82
3944,82
3945,82
3946,82
3947,82
3948,82
3949,82
3950,82
3951,82
3952,82
3953,82
3954,82
3955,82
3956,82
3957,82
3958,82
3959,82
3960,82
3961,82
3962,82
3963,82
3964,82
3965,82
3966,82
3967,82
3968,82
3969,82
3970,82
3971,82
3972,82
3973,82
3974,82
3975,82
3976,82
3977,82
3978,82
3979,82
3980,82
3981,82
3982,82
3983,82
3984,83
3985,83
3986,83
3987,83
3988,83
3989,83
3990,83
3991,83
3992,83
3993,83
3994,83
3995,83
3996,83
3997,83
3998,83
3999,83
4000,83
4001,83
4002,83
4003,83
4004,83
4005,83
4006,83
4007,83
4008,83
4009,83
4010,83
4011,83
4012,83
4013,83
4014,83
4015,83
4016,83
4017,83
4018,83
4019,83
4020,83
4021,83
4022,83
4023,83
4024,83
4025,83
4026,83
4027,83
4028,83
4029,83
4030,83
4031,83
4032,84
4033,84
4034,84
4035,84
4036,84
4037,84
4038,84
4039,84
4040,84
4041,84
4042,84
4043,84
4044,84
4045,84
4046,84
4047,84
4048,84
4049,84
4050,84
4051,84
4052,84
4053,84
4054,84
4055,84
4056,84
4057,84
4058,84
4059,84
4060,84
4061,84
4062,84
4063,84
4064,84
4065,84
4066,84
4067,84
4068,84
4069,84
4070,84
4071,84
4072,84
4073,84
4074,84
4075,84
4076,84
4077,84
4078,84
4079,84
4080,85
4081,85
4082,85
4083,85
4084,85
4085,85
4086,85
4087,85
4088,85
4089,85
4090,85
4091,85
4092,85
4093,85
4094,85
4095,85
4096,85
4097,85
4098,85
4099,85
4100,85
4101,85
4102,85
4103,85
4104,85
4105,85
4106,85
4107,85
4108,85
4109,85
4110,85
4111,85
4112,85
4113,85
4114,85
4115,85
4116,85
4117,85
4118,85
4119,85
4120,85
4121,85
4122,85
4123,85
4124,85
4125,85
4126,85
4127,85
4128,86
4129,86
4130,86
4131,86
4132,86
4133,86
4134,86
4135,86
4136,86
4137,86
4138,86
4139,86
4140,86
4141,86
4142,86
4143,86
4144,86
4145,86
4146,86
4147,86
4148,86
4149,86
4150,86
4151,86
4152,86
4153,86
4154,86
4155,86
4156,86
4157,86
4158,86
4159,86
4160,86
4161,86
4162,86
4163,86
4164,86
4165,86
4166,86
4167,86
4168,86
4169,86
4170,86
4171,86
4172,86
4173,86
4174,86
4175,86
4176,87
4177,87
4178,87
4179,87
4180,87
4181,87
4182,87
4183,87
4184,87
4185,87
4186,87
4187,87
4188,87
4189,87
4190,87
4191,87
4192,87
4193,87
4194,87
4195,87
4196,87
4197,87
4198,87
4199,87
4200,87
4201,87
4202,87
4203,87
4204,87
4205,87
4206,87
4207,87
4208,87
4209,87
4210,87
4211,87
4212,87
4213,87
4214,87
4215,87
4216,87
4217,87
4218,87
4219,87
4220,87
4221,87
4222,87
4223,87
4224,88
4225,88
4226,88
4227,88
4228,88
4229,88
4230,88
4231,88
4232,88
4233,88
4234,88
4235,88
4236,88
4237,88
4238,88
4239,88
4240,88
4241,88
4242,88
4243,88
4244,88
4245,88
4246,88
4247,88
4248,88
4249,88
4250,88
4251,88
4252,88
4253,88
4254,88
4255,88
4256,88
4257,88
4258,88
4259,88
4260,88
4261,88
4262,88
4263,88
4264,88
4265,88
4266,88
4267,88
4268,88
4269,88
4270,88
4271,88
4272,89
4273,89
4274,89
4275,89
4276,89
4277,89
4278,89
4279,89
4280,89
4281,89
4282,89
4283,89
4284,89
4285,89
4286,89
4287,89
4288,89
4289,89
4290,89
4291,89
4292,89
4293,89
4294,89
4295,89
4296,89
4297,89
4298,89
4299,89
4300,89
4301,89
4302,89
4303,89
4304,89
4305,89
4306,89
4307,89
4308,89
4309,89
4310,89
4311,89
4312,89
4313,89
4314,89
4315,89
4316,89
4317,89
4318,89
4319,89
4320,90
4321,90
4322,90
4323,90
4324,90
4325,90
4326,90
4327,90
4328,90
4329,90
4330,90
4331,90
4332,90
4333,90
4334,90
4335,90
4336,90
4337,90
4338,90
4339,90
4340,90
4341,90
4342,90
4343,90
4344,90
4345,90
4346,90
4347,90
4348,90
4349,90
4350,90
4351,90
4352,90
4353,90
4354,90
4355,90
4356,90
4357,90
4358,90
4359,90
4360,90
4361,90
4362,90
4363,90
4364,90
4365,90
4366,90
4367,90
4368,91
4369,91
4370,91
4371,91
4372,91
4373,91
4374,91
4375,91
4376,91
4377,91
4378,91
4379,91
4380,91
4381,91
4382,91
4383,91
4384,91
4385,91
4386,91
4387,91
4388,91
4389,91
4390,91
4391,91
4392,91
4393,91
4394,91
4395,91
4396,91
4397,91
4398,91
4399,91
4400,91
4401,91
4402,91
4403,91
4404,91
4405,91
4406,91
4407,91
4408,91
4409,91
4410,91
4411,91
4412,91
4413,91
4414,91
4415,91
4416,92
4417,92
4418,92
4419,92
4420,92
4421,92
4422,92
4423,92
4424,92
4425,92
4426,92
4427,92
4428,92
4429,92
4430,92
4431,92
4432,92
4433,92
4434,92
4435,92
4436,92
4437,92
4438,92
4439,92
4440,92
4441,92
4442,92
4443,92
4444,92
4445,92
4446,92
4447,92
4448,92
4449,92
4450,92
4451,92
4452,92
4453,92
4454,92
4455,92
4456,92
4457,92
4458,92
4459,92
4460,92
4461,92
4462,92
4463,92
4464,93
4465,93
4466,93
4467,93
4468,93
4469,93
4470,93
4471,93
4472,93
4473,93
4474,93
4475,93
4476,93
4477,93
4478,93
4479,93
4480,93
4481,93
4482,93
4483,93
4484,93
4485,93
4486,93
4487,93
4488,93
4489,93
4490,93
4491,93
4492,93
4493,93
4494,93
4495,93
4496,93
4497,93
4498,93
4499,93
4500,93
4501,93
4502,93
4503,93
4504,93
4505,93
4506,93
4507,93
4508,93
4509,93
4510,93
4511,93
4512,94
4513,94
4514,94
4515,94
4516,94
4517,94
4518,94
4519,94
4520,94
4521,94
4522,94
4523,94
4524,94
4525,94
4526,94
4527,94
4528,94
4529,94
4530,94
4531,94
4532,94
4533,94
4534,94
4535,94
4536,94
4537,94
4538,94
4539,94
4540,94
4541,94
4542,94
4543,94
4544,94
4545,94
4546,94
4547,94
4548,94
4549,94
4550,94
4551,94
4552,94
4553,94
4554,94
4555,94
4556,94
4557,94
4558,94
4559,94
4560,95
4561,95
4562,95
4563,95
4564,95
4565,95
4566,95
4567,95
4568,95
4569,95
4570,95
4571,95
4572,95
4573,95
4574,95
4575,95
4576,95
4577,95
4578,95
4579,95
4580,95
4581,95
4582,95
4583,95
4584,95
4585,95
4586,95
4587,95
4588,95
4589,95
4590,95
4591,95
4592,95
4593,95
4594,95
4595,95
4596,95
4597,95
4598,95
4599,95
4600,95
4601,95
4602,95
4603,95
4604,95
4605,95
4606,95
4607,95
4608,96
4609,96
4610,96
4611,96
4612,96
4613,96
4614,96
4615,96
4616,96
4617,96
4618,96
4619,96
4620,96
4621,96
4622,96
4623,96
4624,96
4625,96
4626,96
4627,96
4628,96
4629,96
4630,96
4631,96
4632,96
4633,96
4634,96
4635,96
4636,96
4637,96
4638,96
4639,96
4640,96
4641,96
4642,96
4643,96
4644,96
4645,96
4646,96
4647,96
4648,96
4649,96
4650,96
4651,96
4652,96
4653,96
4654,96
4655,96
4656,97
4657,97
4658,97
4659,97
4660,97
4661,97
4662,97
4663,97
4664,97
4665,97
4666,97
4667,97
4668,97
4669,97
4670,97
4671,97
4672,97
4673,97
4674,97
4675,97
4676,97
4677,97
4678,97
4679,97
4680,97
4681,97
4682,97
4683,97
4684,97
4685,97
4686,97
4687,97
4688,97
4689,97
4690,97
4691,97
4692,97
4693,97
4694,97
4695,97
4696,97
4697,97
4698,97
4699,97
4700,97
4701,97
4702,97
4703,97
4704,98
4705,98
4706,98
4707,98
4708,98
4709,98
4710,98
4711,98
4712,98
4713,98
4714,98
4715,98
4716,98
4717,98
4718,98
4719,98
4720,98
4721,98
4722,98
4723,98
4724,98
4725,98
4726,98
4727,98
4728,98
4729,98
4730,98
4731,98
4732,98
4733,98
4734,98
4735,98
4736,98
4737,98
4738,98
4739,98
4740,98
4741,98
4742,98
4743,98
4744,98
4745,98
4746,98
4747,98
4748,98
4749,98
4750,98
4751,98
4752,99
4753,99
4754,99
4755,99
4756,99
4757,99
4758,99
4759,99
4760,99
4761,99
4762,99
4763,99
4764,99
4765,99
4766,99
4767,99
4768,99
4769,99
4770,99
4771,99
4772,99
4773,99
4774,99
4775,99
4776,99
4777,99
4778,99
4779,99
4780,99
4781,99
4782,99
4783,99
4784,99
4785,99
4786,99
4787,99
4788,99
4789,99
4790,99
4791,99
4792,99
4793,99
4794,99
4795,99
4796,99
4797,99
4798,99
4799,99
