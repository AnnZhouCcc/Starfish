0,0
1,0
2,0
3,0
4,0
5,0
6,0
7,0
8,0
9,0
10,0
11,0
12,0
13,0
14,0
15,0
16,0
17,0
18,1
19,1
20,1
21,1
22,1
23,1
24,1
25,1
26,1
27,1
28,1
29,1
30,1
31,1
32,1
33,1
34,1
35,1
36,2
37,2
38,2
39,2
40,2
41,2
42,2
43,2
44,2
45,2
46,2
47,2
48,2
49,2
50,2
51,2
52,2
53,2
54,3
55,3
56,3
57,3
58,3
59,3
60,3
61,3
62,3
63,3
64,3
65,3
66,3
67,3
68,3
69,3
70,3
71,3
72,4
73,4
74,4
75,4
76,4
77,4
78,4
79,4
80,4
81,4
82,4
83,4
84,4
85,4
86,4
87,4
88,4
89,4
90,5
91,5
92,5
93,5
94,5
95,5
96,5
97,5
98,5
99,5
100,5
101,5
102,5
103,5
104,5
105,5
106,5
107,5
108,6
109,6
110,6
111,6
112,6
113,6
114,6
115,6
116,6
117,6
118,6
119,6
120,6
121,6
122,6
123,6
124,6
125,6
126,6
127,6
128,7
129,7
130,7
131,7
132,7
133,7
134,7
135,7
136,7
137,7
138,7
139,7
140,7
141,7
142,7
143,7
144,7
145,7
146,7
147,7
148,8
149,8
150,8
151,8
152,8
153,8
154,8
155,8
156,8
157,8
158,8
159,8
160,8
161,8
162,8
163,8
164,8
165,8
166,8
167,8
168,9
169,9
170,9
171,9
172,9
173,9
174,9
175,9
176,9
177,9
178,9
179,9
180,9
181,9
182,9
183,9
184,9
185,9
186,9
187,9
188,10
189,10
190,10
191,10
192,10
193,10
194,10
195,10
196,10
197,10
198,10
199,10
200,10
201,10
202,10
203,10
204,10
205,10
206,11
207,11
208,11
209,11
210,11
211,11
212,11
213,11
214,11
215,11
216,11
217,11
218,11
219,11
220,11
221,11
222,11
223,11
224,12
225,12
226,12
227,12
228,12
229,12
230,12
231,12
232,12
233,12
234,12
235,12
236,12
237,12
238,12
239,12
240,12
241,12
242,13
243,13
244,13
245,13
246,13
247,13
248,13
249,13
250,13
251,13
252,13
253,13
254,13
255,13
256,13
257,13
258,13
259,13
260,14
261,14
262,14
263,14
264,14
265,14
266,14
267,14
268,14
269,14
270,14
271,14
272,14
273,14
274,14
275,14
276,14
277,14
278,15
279,15
280,15
281,15
282,15
283,15
284,15
285,15
286,15
287,15
288,15
289,15
290,15
291,15
292,15
293,15
294,15
295,15
296,16
297,16
298,16
299,16
300,16
301,16
302,16
303,16
304,16
305,16
306,16
307,16
308,16
309,16
310,16
311,16
312,16
313,16
314,16
315,16
316,17
317,17
318,17
319,17
320,17
321,17
322,17
323,17
324,17
325,17
326,17
327,17
328,17
329,17
330,17
331,17
332,17
333,17
334,17
335,17
336,18
337,18
338,18
339,18
340,18
341,18
342,18
343,18
344,18
345,18
346,18
347,18
348,18
349,18
350,18
351,18
352,18
353,18
354,18
355,18
356,19
357,19
358,19
359,19
360,19
361,19
362,19
363,19
364,19
365,19
366,19
367,19
368,19
369,19
370,19
371,19
372,19
373,19
374,19
375,19
376,20
377,20
378,20
379,20
380,20
381,20
382,20
383,20
384,20
385,20
386,20
387,20
388,20
389,20
390,20
391,20
392,20
393,20
394,21
395,21
396,21
397,21
398,21
399,21
400,21
401,21
402,21
403,21
404,21
405,21
406,21
407,21
408,21
409,21
410,21
411,21
412,22
413,22
414,22
415,22
416,22
417,22
418,22
419,22
420,22
421,22
422,22
423,22
424,22
425,22
426,22
427,22
428,22
429,22
430,23
431,23
432,23
433,23
434,23
435,23
436,23
437,23
438,23
439,23
440,23
441,23
442,23
443,23
444,23
445,23
446,23
447,23
448,24
449,24
450,24
451,24
452,24
453,24
454,24
455,24
456,24
457,24
458,24
459,24
460,24
461,24
462,24
463,24
464,24
465,24
466,25
467,25
468,25
469,25
470,25
471,25
472,25
473,25
474,25
475,25
476,25
477,25
478,25
479,25
480,25
481,25
482,25
483,25
484,26
485,26
486,26
487,26
488,26
489,26
490,26
491,26
492,26
493,26
494,26
495,26
496,26
497,26
498,26
499,26
500,26
501,26
502,26
503,26
504,27
505,27
506,27
507,27
508,27
509,27
510,27
511,27
512,27
513,27
514,27
515,27
516,27
517,27
518,27
519,27
520,27
521,27
522,27
523,27
524,28
525,28
526,28
527,28
528,28
529,28
530,28
531,28
532,28
533,28
534,28
535,28
536,28
537,28
538,28
539,28
540,28
541,28
542,28
543,28
544,29
545,29
546,29
547,29
548,29
549,29
550,29
551,29
552,29
553,29
554,29
555,29
556,29
557,29
558,29
559,29
560,29
561,29
562,29
563,29
564,30
565,30
566,30
567,30
568,30
569,30
570,30
571,30
572,30
573,30
574,30
575,30
576,30
577,30
578,30
579,30
580,30
581,30
582,31
583,31
584,31
585,31
586,31
587,31
588,31
589,31
590,31
591,31
592,31
593,31
594,31
595,31
596,31
597,31
598,31
599,31
600,32
601,32
602,32
603,32
604,32
605,32
606,32
607,32
608,32
609,32
610,32
611,32
612,32
613,32
614,32
615,32
616,32
617,32
618,33
619,33
620,33
621,33
622,33
623,33
624,33
625,33
626,33
627,33
628,33
629,33
630,33
631,33
632,33
633,33
634,33
635,33
636,34
637,34
638,34
639,34
640,34
641,34
642,34
643,34
644,34
645,34
646,34
647,34
648,34
649,34
650,34
651,34
652,34
653,34
654,35
655,35
656,35
657,35
658,35
659,35
660,35
661,35
662,35
663,35
664,35
665,35
666,35
667,35
668,35
669,35
670,35
671,35
672,36
673,36
674,36
675,36
676,36
677,36
678,36
679,36
680,36
681,36
682,36
683,36
684,36
685,36
686,36
687,36
688,36
689,36
690,36
691,36
692,37
693,37
694,37
695,37
696,37
697,37
698,37
699,37
700,37
701,37
702,37
703,37
704,37
705,37
706,37
707,37
708,37
709,37
710,37
711,37
712,38
713,38
714,38
715,38
716,38
717,38
718,38
719,38
720,38
721,38
722,38
723,38
724,38
725,38
726,38
727,38
728,38
729,38
730,38
731,38
732,39
733,39
734,39
735,39
736,39
737,39
738,39
739,39
740,39
741,39
742,39
743,39
744,39
745,39
746,39
747,39
748,39
749,39
750,39
751,39
