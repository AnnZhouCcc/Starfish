0,0
1,0
2,0
3,0
4,0
5,0
6,0
7,0
8,0
9,0
10,0
11,0
12,0
13,0
14,0
15,0
16,0
17,0
18,0
19,0
20,0
21,0
22,0
23,0
24,0
25,0
26,0
27,0
28,0
29,0
30,0
31,0
32,0
33,0
34,0
35,0
36,0
37,0
38,0
39,0
40,0
41,0
42,0
43,0
44,0
45,0
46,0
47,0
48,0
49,0
50,0
51,0
52,0
53,0
54,0
55,0
56,1
57,1
58,1
59,1
60,1
61,1
62,1
63,1
64,1
65,1
66,1
67,1
68,1
69,1
70,1
71,1
72,1
73,1
74,1
75,1
76,1
77,1
78,1
79,1
80,1
81,1
82,1
83,1
84,1
85,1
86,1
87,1
88,1
89,1
90,1
91,1
92,1
93,1
94,1
95,1
96,1
97,1
98,1
99,1
100,1
101,1
102,1
103,1
104,1
105,1
106,1
107,1
108,1
109,1
110,1
111,1
112,2
113,2
114,2
115,2
116,2
117,2
118,2
119,2
120,2
121,2
122,2
123,2
124,2
125,2
126,2
127,2
128,2
129,2
130,2
131,2
132,2
133,2
134,2
135,2
136,2
137,2
138,2
139,2
140,2
141,2
142,2
143,2
144,2
145,2
146,2
147,2
148,2
149,2
150,2
151,2
152,2
153,2
154,2
155,2
156,2
157,2
158,2
159,2
160,2
161,2
162,2
163,2
164,2
165,2
166,2
167,2
168,3
169,3
170,3
171,3
172,3
173,3
174,3
175,3
176,3
177,3
178,3
179,3
180,3
181,3
182,3
183,3
184,3
185,3
186,3
187,3
188,3
189,3
190,3
191,3
192,3
193,3
194,3
195,3
196,3
197,3
198,3
199,3
200,3
201,3
202,3
203,3
204,3
205,3
206,3
207,3
208,3
209,3
210,3
211,3
212,3
213,3
214,3
215,3
216,3
217,3
218,3
219,3
220,3
221,3
222,3
223,3
224,4
225,4
226,4
227,4
228,4
229,4
230,4
231,4
232,4
233,4
234,4
235,4
236,4
237,4
238,4
239,4
240,4
241,4
242,4
243,4
244,4
245,4
246,4
247,4
248,4
249,4
250,4
251,4
252,4
253,4
254,4
255,4
256,4
257,4
258,4
259,4
260,4
261,4
262,4
263,4
264,4
265,4
266,4
267,4
268,4
269,4
270,4
271,4
272,4
273,4
274,4
275,4
276,4
277,4
278,4
279,4
280,5
281,5
282,5
283,5
284,5
285,5
286,5
287,5
288,5
289,5
290,5
291,5
292,5
293,5
294,5
295,5
296,5
297,5
298,5
299,5
300,5
301,5
302,5
303,5
304,5
305,5
306,5
307,5
308,5
309,5
310,5
311,5
312,5
313,5
314,5
315,5
316,5
317,5
318,5
319,5
320,5
321,5
322,5
323,5
324,5
325,5
326,5
327,5
328,5
329,5
330,5
331,5
332,5
333,5
334,5
335,5
336,6
337,6
338,6
339,6
340,6
341,6
342,6
343,6
344,6
345,6
346,6
347,6
348,6
349,6
350,6
351,6
352,6
353,6
354,6
355,6
356,6
357,6
358,6
359,6
360,6
361,6
362,6
363,6
364,6
365,6
366,6
367,6
368,6
369,6
370,6
371,6
372,6
373,6
374,6
375,6
376,6
377,6
378,6
379,6
380,6
381,6
382,6
383,6
384,6
385,6
386,6
387,6
388,6
389,6
390,6
391,6
392,7
393,7
394,7
395,7
396,7
397,7
398,7
399,7
400,7
401,7
402,7
403,7
404,7
405,7
406,7
407,7
408,7
409,7
410,7
411,7
412,7
413,7
414,7
415,7
416,7
417,7
418,7
419,7
420,7
421,7
422,7
423,7
424,7
425,7
426,7
427,7
428,7
429,7
430,7
431,7
432,7
433,7
434,7
435,7
436,7
437,7
438,7
439,7
440,7
441,7
442,7
443,7
444,7
445,7
446,7
447,7
448,8
449,8
450,8
451,8
452,8
453,8
454,8
455,8
456,8
457,8
458,8
459,8
460,8
461,8
462,8
463,8
464,8
465,8
466,8
467,8
468,8
469,8
470,8
471,8
472,8
473,8
474,8
475,8
476,8
477,8
478,8
479,8
480,8
481,8
482,8
483,8
484,8
485,8
486,8
487,8
488,8
489,8
490,8
491,8
492,8
493,8
494,8
495,8
496,8
497,8
498,8
499,8
500,8
501,8
502,8
503,8
504,9
505,9
506,9
507,9
508,9
509,9
510,9
511,9
512,9
513,9
514,9
515,9
516,9
517,9
518,9
519,9
520,9
521,9
522,9
523,9
524,9
525,9
526,9
527,9
528,9
529,9
530,9
531,9
532,9
533,9
534,9
535,9
536,9
537,9
538,9
539,9
540,9
541,9
542,9
543,9
544,9
545,9
546,9
547,9
548,9
549,9
550,9
551,9
552,9
553,9
554,9
555,9
556,9
557,9
558,9
559,9
560,10
561,10
562,10
563,10
564,10
565,10
566,10
567,10
568,10
569,10
570,10
571,10
572,10
573,10
574,10
575,10
576,10
577,10
578,10
579,10
580,10
581,10
582,10
583,10
584,10
585,10
586,10
587,10
588,10
589,10
590,10
591,10
592,10
593,10
594,10
595,10
596,10
597,10
598,10
599,10
600,10
601,10
602,10
603,10
604,10
605,10
606,10
607,10
608,10
609,10
610,10
611,10
612,10
613,10
614,10
615,10
616,11
617,11
618,11
619,11
620,11
621,11
622,11
623,11
624,11
625,11
626,11
627,11
628,11
629,11
630,11
631,11
632,11
633,11
634,11
635,11
636,11
637,11
638,11
639,11
640,11
641,11
642,11
643,11
644,11
645,11
646,11
647,11
648,11
649,11
650,11
651,11
652,11
653,11
654,11
655,11
656,11
657,11
658,11
659,11
660,11
661,11
662,11
663,11
664,11
665,11
666,11
667,11
668,11
669,11
670,11
671,11
672,12
673,12
674,12
675,12
676,12
677,12
678,12
679,12
680,12
681,12
682,12
683,12
684,12
685,12
686,12
687,12
688,12
689,12
690,12
691,12
692,12
693,12
694,12
695,12
696,12
697,12
698,12
699,12
700,12
701,12
702,12
703,12
704,12
705,12
706,12
707,12
708,12
709,12
710,12
711,12
712,12
713,12
714,12
715,12
716,12
717,12
718,12
719,12
720,12
721,12
722,12
723,12
724,12
725,12
726,12
727,12
728,13
729,13
730,13
731,13
732,13
733,13
734,13
735,13
736,13
737,13
738,13
739,13
740,13
741,13
742,13
743,13
744,13
745,13
746,13
747,13
748,13
749,13
750,13
751,13
752,13
753,13
754,13
755,13
756,13
757,13
758,13
759,13
760,13
761,13
762,13
763,13
764,13
765,13
766,13
767,13
768,13
769,13
770,13
771,13
772,13
773,13
774,13
775,13
776,13
777,13
778,13
779,13
780,13
781,13
782,13
783,13
784,14
785,14
786,14
787,14
788,14
789,14
790,14
791,14
792,14
793,14
794,14
795,14
796,14
797,14
798,14
799,14
800,14
801,14
802,14
803,14
804,14
805,14
806,14
807,14
808,14
809,14
810,14
811,14
812,14
813,14
814,14
815,14
816,14
817,14
818,14
819,14
820,14
821,14
822,14
823,14
824,14
825,14
826,14
827,14
828,14
829,14
830,14
831,14
832,14
833,14
834,14
835,14
836,14
837,14
838,14
839,14
840,15
841,15
842,15
843,15
844,15
845,15
846,15
847,15
848,15
849,15
850,15
851,15
852,15
853,15
854,15
855,15
856,15
857,15
858,15
859,15
860,15
861,15
862,15
863,15
864,15
865,15
866,15
867,15
868,15
869,15
870,15
871,15
872,15
873,15
874,15
875,15
876,15
877,15
878,15
879,15
880,15
881,15
882,15
883,15
884,15
885,15
886,15
887,15
888,15
889,15
890,15
891,15
892,15
893,15
894,15
895,15
896,16
897,16
898,16
899,16
900,16
901,16
902,16
903,16
904,16
905,16
906,16
907,16
908,16
909,16
910,16
911,16
912,16
913,16
914,16
915,16
916,16
917,16
918,16
919,16
920,16
921,16
922,16
923,16
924,16
925,16
926,16
927,16
928,16
929,16
930,16
931,16
932,16
933,16
934,16
935,16
936,16
937,16
938,16
939,16
940,16
941,16
942,16
943,16
944,16
945,16
946,16
947,16
948,16
949,16
950,16
951,16
952,17
953,17
954,17
955,17
956,17
957,17
958,17
959,17
960,17
961,17
962,17
963,17
964,17
965,17
966,17
967,17
968,17
969,17
970,17
971,17
972,17
973,17
974,17
975,17
976,17
977,17
978,17
979,17
980,17
981,17
982,17
983,17
984,17
985,17
986,17
987,17
988,17
989,17
990,17
991,17
992,17
993,17
994,17
995,17
996,17
997,17
998,17
999,17
1000,17
1001,17
1002,17
1003,17
1004,17
1005,17
1006,17
1007,17
1008,18
1009,18
1010,18
1011,18
1012,18
1013,18
1014,18
1015,18
1016,18
1017,18
1018,18
1019,18
1020,18
1021,18
1022,18
1023,18
1024,18
1025,18
1026,18
1027,18
1028,18
1029,18
1030,18
1031,18
1032,18
1033,18
1034,18
1035,18
1036,18
1037,18
1038,18
1039,18
1040,18
1041,18
1042,18
1043,18
1044,18
1045,18
1046,18
1047,18
1048,18
1049,18
1050,18
1051,18
1052,18
1053,18
1054,18
1055,18
1056,18
1057,18
1058,18
1059,18
1060,18
1061,18
1062,18
1063,18
1064,19
1065,19
1066,19
1067,19
1068,19
1069,19
1070,19
1071,19
1072,19
1073,19
1074,19
1075,19
1076,19
1077,19
1078,19
1079,19
1080,19
1081,19
1082,19
1083,19
1084,19
1085,19
1086,19
1087,19
1088,19
1089,19
1090,19
1091,19
1092,19
1093,19
1094,19
1095,19
1096,19
1097,19
1098,19
1099,19
1100,19
1101,19
1102,19
1103,19
1104,19
1105,19
1106,19
1107,19
1108,19
1109,19
1110,19
1111,19
1112,19
1113,19
1114,19
1115,19
1116,19
1117,19
1118,19
1119,19
1120,20
1121,20
1122,20
1123,20
1124,20
1125,20
1126,20
1127,20
1128,20
1129,20
1130,20
1131,20
1132,20
1133,20
1134,20
1135,20
1136,20
1137,20
1138,20
1139,20
1140,20
1141,20
1142,20
1143,20
1144,20
1145,20
1146,20
1147,20
1148,20
1149,20
1150,20
1151,20
1152,20
1153,20
1154,20
1155,20
1156,20
1157,20
1158,20
1159,20
1160,20
1161,20
1162,20
1163,20
1164,20
1165,20
1166,20
1167,20
1168,20
1169,20
1170,20
1171,20
1172,20
1173,20
1174,20
1175,20
1176,21
1177,21
1178,21
1179,21
1180,21
1181,21
1182,21
1183,21
1184,21
1185,21
1186,21
1187,21
1188,21
1189,21
1190,21
1191,21
1192,21
1193,21
1194,21
1195,21
1196,21
1197,21
1198,21
1199,21
1200,21
1201,21
1202,21
1203,21
1204,21
1205,21
1206,21
1207,21
1208,21
1209,21
1210,21
1211,21
1212,21
1213,21
1214,21
1215,21
1216,21
1217,21
1218,21
1219,21
1220,21
1221,21
1222,21
1223,21
1224,21
1225,21
1226,21
1227,21
1228,21
1229,21
1230,21
1231,21
1232,22
1233,22
1234,22
1235,22
1236,22
1237,22
1238,22
1239,22
1240,22
1241,22
1242,22
1243,22
1244,22
1245,22
1246,22
1247,22
1248,22
1249,22
1250,22
1251,22
1252,22
1253,22
1254,22
1255,22
1256,22
1257,22
1258,22
1259,22
1260,22
1261,22
1262,22
1263,22
1264,22
1265,22
1266,22
1267,22
1268,22
1269,22
1270,22
1271,22
1272,22
1273,22
1274,22
1275,22
1276,22
1277,22
1278,22
1279,22
1280,22
1281,22
1282,22
1283,22
1284,22
1285,22
1286,22
1287,22
1288,23
1289,23
1290,23
1291,23
1292,23
1293,23
1294,23
1295,23
1296,23
1297,23
1298,23
1299,23
1300,23
1301,23
1302,23
1303,23
1304,23
1305,23
1306,23
1307,23
1308,23
1309,23
1310,23
1311,23
1312,23
1313,23
1314,23
1315,23
1316,23
1317,23
1318,23
1319,23
1320,23
1321,23
1322,23
1323,23
1324,23
1325,23
1326,23
1327,23
1328,23
1329,23
1330,23
1331,23
1332,23
1333,23
1334,23
1335,23
1336,23
1337,23
1338,23
1339,23
1340,23
1341,23
1342,23
1343,23
1344,24
1345,24
1346,24
1347,24
1348,24
1349,24
1350,24
1351,24
1352,24
1353,24
1354,24
1355,24
1356,24
1357,24
1358,24
1359,24
1360,24
1361,24
1362,24
1363,24
1364,24
1365,24
1366,24
1367,24
1368,24
1369,24
1370,24
1371,24
1372,24
1373,24
1374,24
1375,24
1376,24
1377,24
1378,24
1379,24
1380,24
1381,24
1382,24
1383,24
1384,24
1385,24
1386,24
1387,24
1388,24
1389,24
1390,24
1391,24
1392,24
1393,24
1394,24
1395,24
1396,24
1397,24
1398,24
1399,24
1400,25
1401,25
1402,25
1403,25
1404,25
1405,25
1406,25
1407,25
1408,25
1409,25
1410,25
1411,25
1412,25
1413,25
1414,25
1415,25
1416,25
1417,25
1418,25
1419,25
1420,25
1421,25
1422,25
1423,25
1424,25
1425,25
1426,25
1427,25
1428,25
1429,25
1430,25
1431,25
1432,25
1433,25
1434,25
1435,25
1436,25
1437,25
1438,25
1439,25
1440,25
1441,25
1442,25
1443,25
1444,25
1445,25
1446,25
1447,25
1448,25
1449,25
1450,25
1451,25
1452,25
1453,25
1454,25
1455,25
1456,26
1457,26
1458,26
1459,26
1460,26
1461,26
1462,26
1463,26
1464,26
1465,26
1466,26
1467,26
1468,26
1469,26
1470,26
1471,26
1472,26
1473,26
1474,26
1475,26
1476,26
1477,26
1478,26
1479,26
1480,26
1481,26
1482,26
1483,26
1484,26
1485,26
1486,26
1487,26
1488,26
1489,26
1490,26
1491,26
1492,26
1493,26
1494,26
1495,26
1496,26
1497,26
1498,26
1499,26
1500,26
1501,26
1502,26
1503,26
1504,26
1505,26
1506,26
1507,26
1508,26
1509,26
1510,26
1511,26
1512,27
1513,27
1514,27
1515,27
1516,27
1517,27
1518,27
1519,27
1520,27
1521,27
1522,27
1523,27
1524,27
1525,27
1526,27
1527,27
1528,27
1529,27
1530,27
1531,27
1532,27
1533,27
1534,27
1535,27
1536,27
1537,27
1538,27
1539,27
1540,27
1541,27
1542,27
1543,27
1544,27
1545,27
1546,27
1547,27
1548,27
1549,27
1550,27
1551,27
1552,27
1553,27
1554,27
1555,27
1556,27
1557,27
1558,27
1559,27
1560,27
1561,27
1562,27
1563,27
1564,27
1565,27
1566,27
1567,27
1568,28
1569,28
1570,28
1571,28
1572,28
1573,28
1574,28
1575,28
1576,28
1577,28
1578,28
1579,28
1580,28
1581,28
1582,28
1583,28
1584,28
1585,28
1586,28
1587,28
1588,28
1589,28
1590,28
1591,28
1592,28
1593,28
1594,28
1595,28
1596,28
1597,28
1598,28
1599,28
1600,28
1601,28
1602,28
1603,28
1604,28
1605,28
1606,28
1607,28
1608,28
1609,28
1610,28
1611,28
1612,28
1613,28
1614,28
1615,28
1616,28
1617,28
1618,28
1619,28
1620,28
1621,28
1622,28
1623,28
1624,29
1625,29
1626,29
1627,29
1628,29
1629,29
1630,29
1631,29
1632,29
1633,29
1634,29
1635,29
1636,29
1637,29
1638,29
1639,29
1640,29
1641,29
1642,29
1643,29
1644,29
1645,29
1646,29
1647,29
1648,29
1649,29
1650,29
1651,29
1652,29
1653,29
1654,29
1655,29
1656,29
1657,29
1658,29
1659,29
1660,29
1661,29
1662,29
1663,29
1664,29
1665,29
1666,29
1667,29
1668,29
1669,29
1670,29
1671,29
1672,29
1673,29
1674,29
1675,29
1676,29
1677,29
1678,29
1679,29
1680,30
1681,30
1682,30
1683,30
1684,30
1685,30
1686,30
1687,30
1688,30
1689,30
1690,30
1691,30
1692,30
1693,30
1694,30
1695,30
1696,30
1697,30
1698,30
1699,30
1700,30
1701,30
1702,30
1703,30
1704,30
1705,30
1706,30
1707,30
1708,30
1709,30
1710,30
1711,30
1712,30
1713,30
1714,30
1715,30
1716,30
1717,30
1718,30
1719,30
1720,30
1721,30
1722,30
1723,30
1724,30
1725,30
1726,30
1727,30
1728,30
1729,30
1730,30
1731,30
1732,30
1733,30
1734,30
1735,30
1736,31
1737,31
1738,31
1739,31
1740,31
1741,31
1742,31
1743,31
1744,31
1745,31
1746,31
1747,31
1748,31
1749,31
1750,31
1751,31
1752,31
1753,31
1754,31
1755,31
1756,31
1757,31
1758,31
1759,31
1760,31
1761,31
1762,31
1763,31
1764,31
1765,31
1766,31
1767,31
1768,31
1769,31
1770,31
1771,31
1772,31
1773,31
1774,31
1775,31
1776,31
1777,31
1778,31
1779,31
1780,31
1781,31
1782,31
1783,31
1784,31
1785,31
1786,31
1787,31
1788,31
1789,31
1790,31
1791,31
1792,32
1793,32
1794,32
1795,32
1796,32
1797,32
1798,32
1799,32
1800,32
1801,32
1802,32
1803,32
1804,32
1805,32
1806,32
1807,32
1808,32
1809,32
1810,32
1811,32
1812,32
1813,32
1814,32
1815,32
1816,32
1817,32
1818,32
1819,32
1820,32
1821,32
1822,32
1823,32
1824,32
1825,32
1826,32
1827,32
1828,32
1829,32
1830,32
1831,32
1832,32
1833,32
1834,32
1835,32
1836,32
1837,32
1838,32
1839,32
1840,32
1841,32
1842,32
1843,32
1844,32
1845,32
1846,32
1847,32
1848,33
1849,33
1850,33
1851,33
1852,33
1853,33
1854,33
1855,33
1856,33
1857,33
1858,33
1859,33
1860,33
1861,33
1862,33
1863,33
1864,33
1865,33
1866,33
1867,33
1868,33
1869,33
1870,33
1871,33
1872,33
1873,33
1874,33
1875,33
1876,33
1877,33
1878,33
1879,33
1880,33
1881,33
1882,33
1883,33
1884,33
1885,33
1886,33
1887,33
1888,33
1889,33
1890,33
1891,33
1892,33
1893,33
1894,33
1895,33
1896,33
1897,33
1898,33
1899,33
1900,33
1901,33
1902,33
1903,33
1904,34
1905,34
1906,34
1907,34
1908,34
1909,34
1910,34
1911,34
1912,34
1913,34
1914,34
1915,34
1916,34
1917,34
1918,34
1919,34
1920,34
1921,34
1922,34
1923,34
1924,34
1925,34
1926,34
1927,34
1928,34
1929,34
1930,34
1931,34
1932,34
1933,34
1934,34
1935,34
1936,34
1937,34
1938,34
1939,34
1940,34
1941,34
1942,34
1943,34
1944,34
1945,34
1946,34
1947,34
1948,34
1949,34
1950,34
1951,34
1952,34
1953,34
1954,34
1955,34
1956,34
1957,34
1958,34
1959,34
1960,35
1961,35
1962,35
1963,35
1964,35
1965,35
1966,35
1967,35
1968,35
1969,35
1970,35
1971,35
1972,35
1973,35
1974,35
1975,35
1976,35
1977,35
1978,35
1979,35
1980,35
1981,35
1982,35
1983,35
1984,35
1985,35
1986,35
1987,35
1988,35
1989,35
1990,35
1991,35
1992,35
1993,35
1994,35
1995,35
1996,35
1997,35
1998,35
1999,35
2000,35
2001,35
2002,35
2003,35
2004,35
2005,35
2006,35
2007,35
2008,35
2009,35
2010,35
2011,35
2012,35
2013,35
2014,35
2015,35
2016,36
2017,36
2018,36
2019,36
2020,36
2021,36
2022,36
2023,36
2024,36
2025,36
2026,36
2027,36
2028,36
2029,36
2030,36
2031,36
2032,36
2033,36
2034,36
2035,36
2036,36
2037,36
2038,36
2039,36
2040,36
2041,36
2042,36
2043,36
2044,36
2045,36
2046,36
2047,36
2048,36
2049,36
2050,36
2051,36
2052,36
2053,36
2054,36
2055,36
2056,36
2057,36
2058,36
2059,36
2060,36
2061,36
2062,36
2063,36
2064,36
2065,36
2066,36
2067,36
2068,36
2069,36
2070,36
2071,36
2072,37
2073,37
2074,37
2075,37
2076,37
2077,37
2078,37
2079,37
2080,37
2081,37
2082,37
2083,37
2084,37
2085,37
2086,37
2087,37
2088,37
2089,37
2090,37
2091,37
2092,37
2093,37
2094,37
2095,37
2096,37
2097,37
2098,37
2099,37
2100,37
2101,37
2102,37
2103,37
2104,37
2105,37
2106,37
2107,37
2108,37
2109,37
2110,37
2111,37
2112,37
2113,37
2114,37
2115,37
2116,37
2117,37
2118,37
2119,37
2120,37
2121,37
2122,37
2123,37
2124,37
2125,37
2126,37
2127,37
2128,38
2129,38
2130,38
2131,38
2132,38
2133,38
2134,38
2135,38
2136,38
2137,38
2138,38
2139,38
2140,38
2141,38
2142,38
2143,38
2144,38
2145,38
2146,38
2147,38
2148,38
2149,38
2150,38
2151,38
2152,38
2153,38
2154,38
2155,38
2156,38
2157,38
2158,38
2159,38
2160,38
2161,38
2162,38
2163,38
2164,38
2165,38
2166,38
2167,38
2168,38
2169,38
2170,38
2171,38
2172,38
2173,38
2174,38
2175,38
2176,38
2177,38
2178,38
2179,38
2180,38
2181,38
2182,38
2183,38
2184,39
2185,39
2186,39
2187,39
2188,39
2189,39
2190,39
2191,39
2192,39
2193,39
2194,39
2195,39
2196,39
2197,39
2198,39
2199,39
2200,39
2201,39
2202,39
2203,39
2204,39
2205,39
2206,39
2207,39
2208,39
2209,39
2210,39
2211,39
2212,39
2213,39
2214,39
2215,39
2216,39
2217,39
2218,39
2219,39
2220,39
2221,39
2222,39
2223,39
2224,39
2225,39
2226,39
2227,39
2228,39
2229,39
2230,39
2231,39
2232,39
2233,39
2234,39
2235,39
2236,39
2237,39
2238,39
2239,39
2240,40
2241,40
2242,40
2243,40
2244,40
2245,40
2246,40
2247,40
2248,40
2249,40
2250,40
2251,40
2252,40
2253,40
2254,40
2255,40
2256,40
2257,40
2258,40
2259,40
2260,40
2261,40
2262,40
2263,40
2264,40
2265,40
2266,40
2267,40
2268,40
2269,40
2270,40
2271,40
2272,40
2273,40
2274,40
2275,40
2276,40
2277,40
2278,40
2279,40
2280,40
2281,40
2282,40
2283,40
2284,40
2285,40
2286,40
2287,40
2288,40
2289,40
2290,40
2291,40
2292,40
2293,40
2294,40
2295,40
2296,41
2297,41
2298,41
2299,41
2300,41
2301,41
2302,41
2303,41
2304,41
2305,41
2306,41
2307,41
2308,41
2309,41
2310,41
2311,41
2312,41
2313,41
2314,41
2315,41
2316,41
2317,41
2318,41
2319,41
2320,41
2321,41
2322,41
2323,41
2324,41
2325,41
2326,41
2327,41
2328,41
2329,41
2330,41
2331,41
2332,41
2333,41
2334,41
2335,41
2336,41
2337,41
2338,41
2339,41
2340,41
2341,41
2342,41
2343,41
2344,41
2345,41
2346,41
2347,41
2348,41
2349,41
2350,41
2351,41
2352,42
2353,42
2354,42
2355,42
2356,42
2357,42
2358,42
2359,42
2360,42
2361,42
2362,42
2363,42
2364,42
2365,42
2366,42
2367,42
2368,42
2369,42
2370,42
2371,42
2372,42
2373,42
2374,42
2375,42
2376,42
2377,42
2378,42
2379,42
2380,42
2381,42
2382,42
2383,42
2384,42
2385,42
2386,42
2387,42
2388,42
2389,42
2390,42
2391,42
2392,42
2393,42
2394,42
2395,42
2396,42
2397,42
2398,42
2399,42
2400,42
2401,42
2402,42
2403,42
2404,42
2405,42
2406,42
2407,42
2408,43
2409,43
2410,43
2411,43
2412,43
2413,43
2414,43
2415,43
2416,43
2417,43
2418,43
2419,43
2420,43
2421,43
2422,43
2423,43
2424,43
2425,43
2426,43
2427,43
2428,43
2429,43
2430,43
2431,43
2432,43
2433,43
2434,43
2435,43
2436,43
2437,43
2438,43
2439,43
2440,43
2441,43
2442,43
2443,43
2444,43
2445,43
2446,43
2447,43
2448,43
2449,43
2450,43
2451,43
2452,43
2453,43
2454,43
2455,43
2456,43
2457,43
2458,43
2459,43
2460,43
2461,43
2462,43
2463,43
2464,44
2465,44
2466,44
2467,44
2468,44
2469,44
2470,44
2471,44
2472,44
2473,44
2474,44
2475,44
2476,44
2477,44
2478,44
2479,44
2480,44
2481,44
2482,44
2483,44
2484,44
2485,44
2486,44
2487,44
2488,44
2489,44
2490,44
2491,44
2492,44
2493,44
2494,44
2495,44
2496,44
2497,44
2498,44
2499,44
2500,44
2501,44
2502,44
2503,44
2504,44
2505,44
2506,44
2507,44
2508,44
2509,44
2510,44
2511,44
2512,44
2513,44
2514,44
2515,44
2516,44
2517,44
2518,44
2519,44
2520,45
2521,45
2522,45
2523,45
2524,45
2525,45
2526,45
2527,45
2528,45
2529,45
2530,45
2531,45
2532,45
2533,45
2534,45
2535,45
2536,45
2537,45
2538,45
2539,45
2540,45
2541,45
2542,45
2543,45
2544,45
2545,45
2546,45
2547,45
2548,45
2549,45
2550,45
2551,45
2552,45
2553,45
2554,45
2555,45
2556,45
2557,45
2558,45
2559,45
2560,45
2561,45
2562,45
2563,45
2564,45
2565,45
2566,45
2567,45
2568,45
2569,45
2570,45
2571,45
2572,45
2573,45
2574,45
2575,45
2576,46
2577,46
2578,46
2579,46
2580,46
2581,46
2582,46
2583,46
2584,46
2585,46
2586,46
2587,46
2588,46
2589,46
2590,46
2591,46
2592,46
2593,46
2594,46
2595,46
2596,46
2597,46
2598,46
2599,46
2600,46
2601,46
2602,46
2603,46
2604,46
2605,46
2606,46
2607,46
2608,46
2609,46
2610,46
2611,46
2612,46
2613,46
2614,46
2615,46
2616,46
2617,46
2618,46
2619,46
2620,46
2621,46
2622,46
2623,46
2624,46
2625,46
2626,46
2627,46
2628,46
2629,46
2630,46
2631,46
2632,47
2633,47
2634,47
2635,47
2636,47
2637,47
2638,47
2639,47
2640,47
2641,47
2642,47
2643,47
2644,47
2645,47
2646,47
2647,47
2648,47
2649,47
2650,47
2651,47
2652,47
2653,47
2654,47
2655,47
2656,47
2657,47
2658,47
2659,47
2660,47
2661,47
2662,47
2663,47
2664,47
2665,47
2666,47
2667,47
2668,47
2669,47
2670,47
2671,47
2672,47
2673,47
2674,47
2675,47
2676,47
2677,47
2678,47
2679,47
2680,47
2681,47
2682,47
2683,47
2684,47
2685,47
2686,47
2687,47
2688,48
2689,48
2690,48
2691,48
2692,48
2693,48
2694,48
2695,48
2696,48
2697,48
2698,48
2699,48
2700,48
2701,48
2702,48
2703,48
2704,48
2705,48
2706,48
2707,48
2708,48
2709,48
2710,48
2711,48
2712,48
2713,48
2714,48
2715,48
2716,48
2717,48
2718,48
2719,48
2720,48
2721,48
2722,48
2723,48
2724,48
2725,48
2726,48
2727,48
2728,48
2729,48
2730,48
2731,48
2732,48
2733,48
2734,48
2735,48
2736,48
2737,48
2738,48
2739,48
2740,48
2741,48
2742,48
2743,48
2744,49
2745,49
2746,49
2747,49
2748,49
2749,49
2750,49
2751,49
2752,49
2753,49
2754,49
2755,49
2756,49
2757,49
2758,49
2759,49
2760,49
2761,49
2762,49
2763,49
2764,49
2765,49
2766,49
2767,49
2768,49
2769,49
2770,49
2771,49
2772,49
2773,49
2774,49
2775,49
2776,49
2777,49
2778,49
2779,49
2780,49
2781,49
2782,49
2783,49
2784,49
2785,49
2786,49
2787,49
2788,49
2789,49
2790,49
2791,49
2792,49
2793,49
2794,49
2795,49
2796,49
2797,49
2798,49
2799,49
2800,50
2801,50
2802,50
2803,50
2804,50
2805,50
2806,50
2807,50
2808,50
2809,50
2810,50
2811,50
2812,50
2813,50
2814,50
2815,50
2816,50
2817,50
2818,50
2819,50
2820,50
2821,50
2822,50
2823,50
2824,50
2825,50
2826,50
2827,50
2828,50
2829,50
2830,50
2831,50
2832,50
2833,50
2834,50
2835,50
2836,50
2837,50
2838,50
2839,50
2840,50
2841,50
2842,50
2843,50
2844,50
2845,50
2846,50
2847,50
2848,50
2849,50
2850,50
2851,50
2852,50
2853,50
2854,50
2855,50
2856,51
2857,51
2858,51
2859,51
2860,51
2861,51
2862,51
2863,51
2864,51
2865,51
2866,51
2867,51
2868,51
2869,51
2870,51
2871,51
2872,51
2873,51
2874,51
2875,51
2876,51
2877,51
2878,51
2879,51
2880,51
2881,51
2882,51
2883,51
2884,51
2885,51
2886,51
2887,51
2888,51
2889,51
2890,51
2891,51
2892,51
2893,51
2894,51
2895,51
2896,51
2897,51
2898,51
2899,51
2900,51
2901,51
2902,51
2903,51
2904,51
2905,51
2906,51
2907,51
2908,51
2909,51
2910,51
2911,51
2912,52
2913,52
2914,52
2915,52
2916,52
2917,52
2918,52
2919,52
2920,52
2921,52
2922,52
2923,52
2924,52
2925,52
2926,52
2927,52
2928,52
2929,52
2930,52
2931,52
2932,52
2933,52
2934,52
2935,52
2936,52
2937,52
2938,52
2939,52
2940,52
2941,52
2942,52
2943,52
2944,52
2945,52
2946,52
2947,52
2948,52
2949,52
2950,52
2951,52
2952,52
2953,52
2954,52
2955,52
2956,52
2957,52
2958,52
2959,52
2960,52
2961,52
2962,52
2963,52
2964,52
2965,52
2966,52
2967,52
2968,53
2969,53
2970,53
2971,53
2972,53
2973,53
2974,53
2975,53
2976,53
2977,53
2978,53
2979,53
2980,53
2981,53
2982,53
2983,53
2984,53
2985,53
2986,53
2987,53
2988,53
2989,53
2990,53
2991,53
2992,53
2993,53
2994,53
2995,53
2996,53
2997,53
2998,53
2999,53
3000,53
3001,53
3002,53
3003,53
3004,53
3005,53
3006,53
3007,53
3008,53
3009,53
3010,53
3011,53
3012,53
3013,53
3014,53
3015,53
3016,53
3017,53
3018,53
3019,53
3020,53
3021,53
3022,53
3023,53
3024,54
3025,54
3026,54
3027,54
3028,54
3029,54
3030,54
3031,54
3032,54
3033,54
3034,54
3035,54
3036,54
3037,54
3038,54
3039,54
3040,54
3041,54
3042,54
3043,54
3044,54
3045,54
3046,54
3047,54
3048,54
3049,54
3050,54
3051,54
3052,54
3053,54
3054,54
3055,54
3056,54
3057,54
3058,54
3059,54
3060,54
3061,54
3062,54
3063,54
3064,54
3065,54
3066,54
3067,54
3068,54
3069,54
3070,54
3071,54
3072,54
3073,54
3074,54
3075,54
3076,54
3077,54
3078,54
3079,54
3080,55
3081,55
3082,55
3083,55
3084,55
3085,55
3086,55
3087,55
3088,55
3089,55
3090,55
3091,55
3092,55
3093,55
3094,55
3095,55
3096,55
3097,55
3098,55
3099,55
3100,55
3101,55
3102,55
3103,55
3104,55
3105,55
3106,55
3107,55
3108,55
3109,55
3110,55
3111,55
3112,55
3113,55
3114,55
3115,55
3116,55
3117,55
3118,55
3119,55
3120,55
3121,55
3122,55
3123,55
3124,55
3125,55
3126,55
3127,55
3128,55
3129,55
3130,55
3131,55
3132,55
3133,55
3134,55
3135,55
3136,56
3137,56
3138,56
3139,56
3140,56
3141,56
3142,56
3143,56
3144,56
3145,56
3146,56
3147,56
3148,56
3149,56
3150,56
3151,56
3152,56
3153,56
3154,56
3155,56
3156,56
3157,56
3158,56
3159,56
3160,56
3161,56
3162,56
3163,56
3164,56
3165,56
3166,56
3167,56
3168,56
3169,56
3170,56
3171,56
3172,56
3173,56
3174,56
3175,56
3176,56
3177,56
3178,56
3179,56
3180,56
3181,56
3182,56
3183,56
3184,56
3185,56
3186,56
3187,56
3188,56
3189,56
3190,56
3191,56
3192,57
3193,57
3194,57
3195,57
3196,57
3197,57
3198,57
3199,57
3200,57
3201,57
3202,57
3203,57
3204,57
3205,57
3206,57
3207,57
3208,57
3209,57
3210,57
3211,57
3212,57
3213,57
3214,57
3215,57
3216,57
3217,57
3218,57
3219,57
3220,57
3221,57
3222,57
3223,57
3224,57
3225,57
3226,57
3227,57
3228,57
3229,57
3230,57
3231,57
3232,57
3233,57
3234,57
3235,57
3236,57
3237,57
3238,57
3239,57
3240,57
3241,57
3242,57
3243,57
3244,57
3245,57
3246,57
3247,57
3248,58
3249,58
3250,58
3251,58
3252,58
3253,58
3254,58
3255,58
3256,58
3257,58
3258,58
3259,58
3260,58
3261,58
3262,58
3263,58
3264,58
3265,58
3266,58
3267,58
3268,58
3269,58
3270,58
3271,58
3272,58
3273,58
3274,58
3275,58
3276,58
3277,58
3278,58
3279,58
3280,58
3281,58
3282,58
3283,58
3284,58
3285,58
3286,58
3287,58
3288,58
3289,58
3290,58
3291,58
3292,58
3293,58
3294,58
3295,58
3296,58
3297,58
3298,58
3299,58
3300,58
3301,58
3302,58
3303,58
3304,59
3305,59
3306,59
3307,59
3308,59
3309,59
3310,59
3311,59
3312,59
3313,59
3314,59
3315,59
3316,59
3317,59
3318,59
3319,59
3320,59
3321,59
3322,59
3323,59
3324,59
3325,59
3326,59
3327,59
3328,59
3329,59
3330,59
3331,59
3332,59
3333,59
3334,59
3335,59
3336,59
3337,59
3338,59
3339,59
3340,59
3341,59
3342,59
3343,59
3344,59
3345,59
3346,59
3347,59
3348,59
3349,59
3350,59
3351,59
3352,59
3353,59
3354,59
3355,59
3356,59
3357,59
3358,59
3359,59
3360,60
3361,60
3362,60
3363,60
3364,60
3365,60
3366,60
3367,60
3368,60
3369,60
3370,60
3371,60
3372,60
3373,60
3374,60
3375,60
3376,60
3377,60
3378,60
3379,60
3380,60
3381,60
3382,60
3383,60
3384,60
3385,60
3386,60
3387,60
3388,60
3389,60
3390,60
3391,60
3392,60
3393,60
3394,60
3395,60
3396,60
3397,60
3398,60
3399,60
3400,60
3401,60
3402,60
3403,60
3404,60
3405,60
3406,60
3407,60
3408,60
3409,60
3410,60
3411,60
3412,60
3413,60
3414,60
3415,60
3416,61
3417,61
3418,61
3419,61
3420,61
3421,61
3422,61
3423,61
3424,61
3425,61
3426,61
3427,61
3428,61
3429,61
3430,61
3431,61
3432,61
3433,61
3434,61
3435,61
3436,61
3437,61
3438,61
3439,61
3440,61
3441,61
3442,61
3443,61
3444,61
3445,61
3446,61
3447,61
3448,61
3449,61
3450,61
3451,61
3452,61
3453,61
3454,61
3455,61
3456,61
3457,61
3458,61
3459,61
3460,61
3461,61
3462,61
3463,61
3464,61
3465,61
3466,61
3467,61
3468,61
3469,61
3470,61
3471,61
3472,62
3473,62
3474,62
3475,62
3476,62
3477,62
3478,62
3479,62
3480,62
3481,62
3482,62
3483,62
3484,62
3485,62
3486,62
3487,62
3488,62
3489,62
3490,62
3491,62
3492,62
3493,62
3494,62
3495,62
3496,62
3497,62
3498,62
3499,62
3500,62
3501,62
3502,62
3503,62
3504,62
3505,62
3506,62
3507,62
3508,62
3509,62
3510,62
3511,62
3512,62
3513,62
3514,62
3515,62
3516,62
3517,62
3518,62
3519,62
3520,62
3521,62
3522,62
3523,62
3524,62
3525,62
3526,62
3527,62
3528,63
3529,63
3530,63
3531,63
3532,63
3533,63
3534,63
3535,63
3536,63
3537,63
3538,63
3539,63
3540,63
3541,63
3542,63
3543,63
3544,63
3545,63
3546,63
3547,63
3548,63
3549,63
3550,63
3551,63
3552,63
3553,63
3554,63
3555,63
3556,63
3557,63
3558,63
3559,63
3560,63
3561,63
3562,63
3563,63
3564,63
3565,63
3566,63
3567,63
3568,63
3569,63
3570,63
3571,63
3572,63
3573,63
3574,63
3575,63
3576,63
3577,63
3578,63
3579,63
3580,63
3581,63
3582,63
3583,63
3584,64
3585,64
3586,64
3587,64
3588,64
3589,64
3590,64
3591,64
3592,64
3593,64
3594,64
3595,64
3596,64
3597,64
3598,64
3599,64
3600,64
3601,64
3602,64
3603,64
3604,64
3605,64
3606,64
3607,64
3608,64
3609,64
3610,64
3611,64
3612,64
3613,64
3614,64
3615,64
3616,64
3617,64
3618,64
3619,64
3620,64
3621,64
3622,64
3623,64
3624,64
3625,64
3626,64
3627,64
3628,64
3629,64
3630,64
3631,64
3632,64
3633,64
3634,64
3635,64
3636,64
3637,64
3638,64
3639,64
3640,65
3641,65
3642,65
3643,65
3644,65
3645,65
3646,65
3647,65
3648,65
3649,65
3650,65
3651,65
3652,65
3653,65
3654,65
3655,65
3656,65
3657,65
3658,65
3659,65
3660,65
3661,65
3662,65
3663,65
3664,65
3665,65
3666,65
3667,65
3668,65
3669,65
3670,65
3671,65
3672,65
3673,65
3674,65
3675,65
3676,65
3677,65
3678,65
3679,65
3680,65
3681,65
3682,65
3683,65
3684,65
3685,65
3686,65
3687,65
3688,65
3689,65
3690,65
3691,65
3692,65
3693,65
3694,65
3695,65
3696,66
3697,66
3698,66
3699,66
3700,66
3701,66
3702,66
3703,66
3704,66
3705,66
3706,66
3707,66
3708,66
3709,66
3710,66
3711,66
3712,66
3713,66
3714,66
3715,66
3716,66
3717,66
3718,66
3719,66
3720,66
3721,66
3722,66
3723,66
3724,66
3725,66
3726,66
3727,66
3728,66
3729,66
3730,66
3731,66
3732,66
3733,66
3734,66
3735,66
3736,66
3737,66
3738,66
3739,66
3740,66
3741,66
3742,66
3743,66
3744,66
3745,66
3746,66
3747,66
3748,66
3749,66
3750,66
3751,66
3752,67
3753,67
3754,67
3755,67
3756,67
3757,67
3758,67
3759,67
3760,67
3761,67
3762,67
3763,67
3764,67
3765,67
3766,67
3767,67
3768,67
3769,67
3770,67
3771,67
3772,67
3773,67
3774,67
3775,67
3776,67
3777,67
3778,67
3779,67
3780,67
3781,67
3782,67
3783,67
3784,67
3785,67
3786,67
3787,67
3788,67
3789,67
3790,67
3791,67
3792,67
3793,67
3794,67
3795,67
3796,67
3797,67
3798,67
3799,67
3800,67
3801,67
3802,67
3803,67
3804,67
3805,67
3806,67
3807,67
3808,68
3809,68
3810,68
3811,68
3812,68
3813,68
3814,68
3815,68
3816,68
3817,68
3818,68
3819,68
3820,68
3821,68
3822,68
3823,68
3824,68
3825,68
3826,68
3827,68
3828,68
3829,68
3830,68
3831,68
3832,68
3833,68
3834,68
3835,68
3836,68
3837,68
3838,68
3839,68
3840,68
3841,68
3842,68
3843,68
3844,68
3845,68
3846,68
3847,68
3848,68
3849,68
3850,68
3851,68
3852,68
3853,68
3854,68
3855,68
3856,68
3857,68
3858,68
3859,68
3860,68
3861,68
3862,68
3863,68
3864,69
3865,69
3866,69
3867,69
3868,69
3869,69
3870,69
3871,69
3872,69
3873,69
3874,69
3875,69
3876,69
3877,69
3878,69
3879,69
3880,69
3881,69
3882,69
3883,69
3884,69
3885,69
3886,69
3887,69
3888,69
3889,69
3890,69
3891,69
3892,69
3893,69
3894,69
3895,69
3896,69
3897,69
3898,69
3899,69
3900,69
3901,69
3902,69
3903,69
3904,69
3905,69
3906,69
3907,69
3908,69
3909,69
3910,69
3911,69
3912,69
3913,69
3914,69
3915,69
3916,69
3917,69
3918,69
3919,69
3920,70
3921,70
3922,70
3923,70
3924,70
3925,70
3926,70
3927,70
3928,70
3929,70
3930,70
3931,70
3932,70
3933,70
3934,70
3935,70
3936,70
3937,70
3938,70
3939,70
3940,70
3941,70
3942,70
3943,70
3944,70
3945,70
3946,70
3947,70
3948,70
3949,70
3950,70
3951,70
3952,70
3953,70
3954,70
3955,70
3956,70
3957,70
3958,70
3959,70
3960,70
3961,70
3962,70
3963,70
3964,70
3965,70
3966,70
3967,70
3968,70
3969,70
3970,70
3971,70
3972,70
3973,70
3974,70
3975,70
3976,71
3977,71
3978,71
3979,71
3980,71
3981,71
3982,71
3983,71
3984,71
3985,71
3986,71
3987,71
3988,71
3989,71
3990,71
3991,71
3992,71
3993,71
3994,71
3995,71
3996,71
3997,71
3998,71
3999,71
4000,71
4001,71
4002,71
4003,71
4004,71
4005,71
4006,71
4007,71
4008,71
4009,71
4010,71
4011,71
4012,71
4013,71
4014,71
4015,71
4016,71
4017,71
4018,71
4019,71
4020,71
4021,71
4022,71
4023,71
4024,71
4025,71
4026,71
4027,71
4028,71
4029,71
4030,71
4031,71
4032,72
4033,72
4034,72
4035,72
4036,72
4037,72
4038,72
4039,72
4040,72
4041,72
4042,72
4043,72
4044,72
4045,72
4046,72
4047,72
4048,72
4049,72
4050,72
4051,72
4052,72
4053,72
4054,72
4055,72
4056,72
4057,72
4058,72
4059,72
4060,72
4061,72
4062,72
4063,72
4064,72
4065,72
4066,72
4067,72
4068,72
4069,72
4070,72
4071,72
4072,72
4073,72
4074,72
4075,72
4076,72
4077,72
4078,72
4079,72
4080,72
4081,72
4082,72
4083,72
4084,72
4085,72
4086,72
4087,72
4088,73
4089,73
4090,73
4091,73
4092,73
4093,73
4094,73
4095,73
4096,73
4097,73
4098,73
4099,73
4100,73
4101,73
4102,73
4103,73
4104,73
4105,73
4106,73
4107,73
4108,73
4109,73
4110,73
4111,73
4112,73
4113,73
4114,73
4115,73
4116,73
4117,73
4118,73
4119,73
4120,73
4121,73
4122,73
4123,73
4124,73
4125,73
4126,73
4127,73
4128,73
4129,73
4130,73
4131,73
4132,73
4133,73
4134,73
4135,73
4136,73
4137,73
4138,73
4139,73
4140,73
4141,73
4142,73
4143,73
4144,74
4145,74
4146,74
4147,74
4148,74
4149,74
4150,74
4151,74
4152,74
4153,74
4154,74
4155,74
4156,74
4157,74
4158,74
4159,74
4160,74
4161,74
4162,74
4163,74
4164,74
4165,74
4166,74
4167,74
4168,74
4169,74
4170,74
4171,74
4172,74
4173,74
4174,74
4175,74
4176,74
4177,74
4178,74
4179,74
4180,74
4181,74
4182,74
4183,74
4184,74
4185,74
4186,74
4187,74
4188,74
4189,74
4190,74
4191,74
4192,74
4193,74
4194,74
4195,74
4196,74
4197,74
4198,74
4199,74
4200,75
4201,75
4202,75
4203,75
4204,75
4205,75
4206,75
4207,75
4208,75
4209,75
4210,75
4211,75
4212,75
4213,75
4214,75
4215,75
4216,75
4217,75
4218,75
4219,75
4220,75
4221,75
4222,75
4223,75
4224,75
4225,75
4226,75
4227,75
4228,75
4229,75
4230,75
4231,75
4232,75
4233,75
4234,75
4235,75
4236,75
4237,75
4238,75
4239,75
4240,75
4241,75
4242,75
4243,75
4244,75
4245,75
4246,75
4247,75
4248,75
4249,75
4250,75
4251,75
4252,75
4253,75
4254,75
4255,75
4256,76
4257,76
4258,76
4259,76
4260,76
4261,76
4262,76
4263,76
4264,76
4265,76
4266,76
4267,76
4268,76
4269,76
4270,76
4271,76
4272,76
4273,76
4274,76
4275,76
4276,76
4277,76
4278,76
4279,76
4280,76
4281,76
4282,76
4283,76
4284,76
4285,76
4286,76
4287,76
4288,76
4289,76
4290,76
4291,76
4292,76
4293,76
4294,76
4295,76
4296,76
4297,76
4298,76
4299,76
4300,76
4301,76
4302,76
4303,76
4304,76
4305,76
4306,76
4307,76
4308,76
4309,76
4310,76
4311,76
4312,77
4313,77
4314,77
4315,77
4316,77
4317,77
4318,77
4319,77
4320,77
4321,77
4322,77
4323,77
4324,77
4325,77
4326,77
4327,77
4328,77
4329,77
4330,77
4331,77
4332,77
4333,77
4334,77
4335,77
4336,77
4337,77
4338,77
4339,77
4340,77
4341,77
4342,77
4343,77
4344,77
4345,77
4346,77
4347,77
4348,77
4349,77
4350,77
4351,77
4352,77
4353,77
4354,77
4355,77
4356,77
4357,77
4358,77
4359,77
4360,77
4361,77
4362,77
4363,77
4364,77
4365,77
4366,77
4367,77
4368,78
4369,78
4370,78
4371,78
4372,78
4373,78
4374,78
4375,78
4376,78
4377,78
4378,78
4379,78
4380,78
4381,78
4382,78
4383,78
4384,78
4385,78
4386,78
4387,78
4388,78
4389,78
4390,78
4391,78
4392,78
4393,78
4394,78
4395,78
4396,78
4397,78
4398,78
4399,78
4400,78
4401,78
4402,78
4403,78
4404,78
4405,78
4406,78
4407,78
4408,78
4409,78
4410,78
4411,78
4412,78
4413,78
4414,78
4415,78
4416,78
4417,78
4418,78
4419,78
4420,78
4421,78
4422,78
4423,78
4424,79
4425,79
4426,79
4427,79
4428,79
4429,79
4430,79
4431,79
4432,79
4433,79
4434,79
4435,79
4436,79
4437,79
4438,79
4439,79
4440,79
4441,79
4442,79
4443,79
4444,79
4445,79
4446,79
4447,79
4448,79
4449,79
4450,79
4451,79
4452,79
4453,79
4454,79
4455,79
4456,79
4457,79
4458,79
4459,79
4460,79
4461,79
4462,79
4463,79
4464,79
4465,79
4466,79
4467,79
4468,79
4469,79
4470,79
4471,79
4472,79
4473,79
4474,79
4475,79
4476,79
4477,79
4478,79
4479,79
4480,80
4481,80
4482,80
4483,80
4484,80
4485,80
4486,80
4487,80
4488,80
4489,80
4490,80
4491,80
4492,80
4493,80
4494,80
4495,80
4496,80
4497,80
4498,80
4499,80
4500,80
4501,80
4502,80
4503,80
4504,80
4505,80
4506,80
4507,80
4508,80
4509,80
4510,80
4511,80
4512,80
4513,80
4514,80
4515,80
4516,80
4517,80
4518,80
4519,80
4520,80
4521,80
4522,80
4523,80
4524,80
4525,80
4526,80
4527,80
4528,80
4529,80
4530,80
4531,80
4532,80
4533,80
4534,80
4535,80
4536,81
4537,81
4538,81
4539,81
4540,81
4541,81
4542,81
4543,81
4544,81
4545,81
4546,81
4547,81
4548,81
4549,81
4550,81
4551,81
4552,81
4553,81
4554,81
4555,81
4556,81
4557,81
4558,81
4559,81
4560,81
4561,81
4562,81
4563,81
4564,81
4565,81
4566,81
4567,81
4568,81
4569,81
4570,81
4571,81
4572,81
4573,81
4574,81
4575,81
4576,81
4577,81
4578,81
4579,81
4580,81
4581,81
4582,81
4583,81
4584,81
4585,81
4586,81
4587,81
4588,81
4589,81
4590,81
4591,81
4592,82
4593,82
4594,82
4595,82
4596,82
4597,82
4598,82
4599,82
4600,82
4601,82
4602,82
4603,82
4604,82
4605,82
4606,82
4607,82
4608,82
4609,82
4610,82
4611,82
4612,82
4613,82
4614,82
4615,82
4616,82
4617,82
4618,82
4619,82
4620,82
4621,82
4622,82
4623,82
4624,82
4625,82
4626,82
4627,82
4628,82
4629,82
4630,82
4631,82
4632,82
4633,82
4634,82
4635,82
4636,82
4637,82
4638,82
4639,82
4640,82
4641,82
4642,82
4643,82
4644,82
4645,82
4646,82
4647,82
4648,83
4649,83
4650,83
4651,83
4652,83
4653,83
4654,83
4655,83
4656,83
4657,83
4658,83
4659,83
4660,83
4661,83
4662,83
4663,83
4664,83
4665,83
4666,83
4667,83
4668,83
4669,83
4670,83
4671,83
4672,83
4673,83
4674,83
4675,83
4676,83
4677,83
4678,83
4679,83
4680,83
4681,83
4682,83
4683,83
4684,83
4685,83
4686,83
4687,83
4688,83
4689,83
4690,83
4691,83
4692,83
4693,83
4694,83
4695,83
4696,83
4697,83
4698,83
4699,83
4700,83
4701,83
4702,83
4703,83
4704,84
4705,84
4706,84
4707,84
4708,84
4709,84
4710,84
4711,84
4712,84
4713,84
4714,84
4715,84
4716,84
4717,84
4718,84
4719,84
4720,84
4721,84
4722,84
4723,84
4724,84
4725,84
4726,84
4727,84
4728,84
4729,84
4730,84
4731,84
4732,84
4733,84
4734,84
4735,84
4736,84
4737,84
4738,84
4739,84
4740,84
4741,84
4742,84
4743,84
4744,84
4745,84
4746,84
4747,84
4748,84
4749,84
4750,84
4751,84
4752,84
4753,84
4754,84
4755,84
4756,84
4757,84
4758,84
4759,84
4760,85
4761,85
4762,85
4763,85
4764,85
4765,85
4766,85
4767,85
4768,85
4769,85
4770,85
4771,85
4772,85
4773,85
4774,85
4775,85
4776,85
4777,85
4778,85
4779,85
4780,85
4781,85
4782,85
4783,85
4784,85
4785,85
4786,85
4787,85
4788,85
4789,85
4790,85
4791,85
4792,85
4793,85
4794,85
4795,85
4796,85
4797,85
4798,85
4799,85
4800,85
4801,85
4802,85
4803,85
4804,85
4805,85
4806,85
4807,85
4808,85
4809,85
4810,85
4811,85
4812,85
4813,85
4814,85
4815,85
4816,86
4817,86
4818,86
4819,86
4820,86
4821,86
4822,86
4823,86
4824,86
4825,86
4826,86
4827,86
4828,86
4829,86
4830,86
4831,86
4832,86
4833,86
4834,86
4835,86
4836,86
4837,86
4838,86
4839,86
4840,86
4841,86
4842,86
4843,86
4844,86
4845,86
4846,86
4847,86
4848,86
4849,86
4850,86
4851,86
4852,86
4853,86
4854,86
4855,86
4856,86
4857,86
4858,86
4859,86
4860,86
4861,86
4862,86
4863,86
4864,86
4865,86
4866,86
4867,86
4868,86
4869,86
4870,86
4871,86
4872,87
4873,87
4874,87
4875,87
4876,87
4877,87
4878,87
4879,87
4880,87
4881,87
4882,87
4883,87
4884,87
4885,87
4886,87
4887,87
4888,87
4889,87
4890,87
4891,87
4892,87
4893,87
4894,87
4895,87
4896,87
4897,87
4898,87
4899,87
4900,87
4901,87
4902,87
4903,87
4904,87
4905,87
4906,87
4907,87
4908,87
4909,87
4910,87
4911,87
4912,87
4913,87
4914,87
4915,87
4916,87
4917,87
4918,87
4919,87
4920,87
4921,87
4922,87
4923,87
4924,87
4925,87
4926,87
4927,87
4928,88
4929,88
4930,88
4931,88
4932,88
4933,88
4934,88
4935,88
4936,88
4937,88
4938,88
4939,88
4940,88
4941,88
4942,88
4943,88
4944,88
4945,88
4946,88
4947,88
4948,88
4949,88
4950,88
4951,88
4952,88
4953,88
4954,88
4955,88
4956,88
4957,88
4958,88
4959,88
4960,88
4961,88
4962,88
4963,88
4964,88
4965,88
4966,88
4967,88
4968,88
4969,88
4970,88
4971,88
4972,88
4973,88
4974,88
4975,88
4976,88
4977,88
4978,88
4979,88
4980,88
4981,88
4982,88
4983,88
4984,89
4985,89
4986,89
4987,89
4988,89
4989,89
4990,89
4991,89
4992,89
4993,89
4994,89
4995,89
4996,89
4997,89
4998,89
4999,89
5000,89
5001,89
5002,89
5003,89
5004,89
5005,89
5006,89
5007,89
5008,89
5009,89
5010,89
5011,89
5012,89
5013,89
5014,89
5015,89
5016,89
5017,89
5018,89
5019,89
5020,89
5021,89
5022,89
5023,89
5024,89
5025,89
5026,89
5027,89
5028,89
5029,89
5030,89
5031,89
5032,89
5033,89
5034,89
5035,89
5036,89
5037,89
5038,89
5039,89
5040,90
5041,90
5042,90
5043,90
5044,90
5045,90
5046,90
5047,90
5048,90
5049,90
5050,90
5051,90
5052,90
5053,90
5054,90
5055,90
5056,90
5057,90
5058,90
5059,90
5060,90
5061,90
5062,90
5063,90
5064,90
5065,90
5066,90
5067,90
5068,90
5069,90
5070,90
5071,90
5072,90
5073,90
5074,90
5075,90
5076,90
5077,90
5078,90
5079,90
5080,90
5081,90
5082,90
5083,90
5084,90
5085,90
5086,90
5087,90
5088,90
5089,90
5090,90
5091,90
5092,90
5093,90
5094,90
5095,90
5096,91
5097,91
5098,91
5099,91
5100,91
5101,91
5102,91
5103,91
5104,91
5105,91
5106,91
5107,91
5108,91
5109,91
5110,91
5111,91
5112,91
5113,91
5114,91
5115,91
5116,91
5117,91
5118,91
5119,91
5120,91
5121,91
5122,91
5123,91
5124,91
5125,91
5126,91
5127,91
5128,91
5129,91
5130,91
5131,91
5132,91
5133,91
5134,91
5135,91
5136,91
5137,91
5138,91
5139,91
5140,91
5141,91
5142,91
5143,91
5144,91
5145,91
5146,91
5147,91
5148,91
5149,91
5150,91
5151,91
5152,92
5153,92
5154,92
5155,92
5156,92
5157,92
5158,92
5159,92
5160,92
5161,92
5162,92
5163,92
5164,92
5165,92
5166,92
5167,92
5168,92
5169,92
5170,92
5171,92
5172,92
5173,92
5174,92
5175,92
5176,92
5177,92
5178,92
5179,92
5180,92
5181,92
5182,92
5183,92
5184,92
5185,92
5186,92
5187,92
5188,92
5189,92
5190,92
5191,92
5192,92
5193,92
5194,92
5195,92
5196,92
5197,92
5198,92
5199,92
5200,92
5201,92
5202,92
5203,92
5204,92
5205,92
5206,92
5207,92
5208,93
5209,93
5210,93
5211,93
5212,93
5213,93
5214,93
5215,93
5216,93
5217,93
5218,93
5219,93
5220,93
5221,93
5222,93
5223,93
5224,93
5225,93
5226,93
5227,93
5228,93
5229,93
5230,93
5231,93
5232,93
5233,93
5234,93
5235,93
5236,93
5237,93
5238,93
5239,93
5240,93
5241,93
5242,93
5243,93
5244,93
5245,93
5246,93
5247,93
5248,93
5249,93
5250,93
5251,93
5252,93
5253,93
5254,93
5255,93
5256,93
5257,93
5258,93
5259,93
5260,93
5261,93
5262,93
5263,93
5264,94
5265,94
5266,94
5267,94
5268,94
5269,94
5270,94
5271,94
5272,94
5273,94
5274,94
5275,94
5276,94
5277,94
5278,94
5279,94
5280,94
5281,94
5282,94
5283,94
5284,94
5285,94
5286,94
5287,94
5288,94
5289,94
5290,94
5291,94
5292,94
5293,94
5294,94
5295,94
5296,94
5297,94
5298,94
5299,94
5300,94
5301,94
5302,94
5303,94
5304,94
5305,94
5306,94
5307,94
5308,94
5309,94
5310,94
5311,94
5312,94
5313,94
5314,94
5315,94
5316,94
5317,94
5318,94
5319,94
5320,95
5321,95
5322,95
5323,95
5324,95
5325,95
5326,95
5327,95
5328,95
5329,95
5330,95
5331,95
5332,95
5333,95
5334,95
5335,95
5336,95
5337,95
5338,95
5339,95
5340,95
5341,95
5342,95
5343,95
5344,95
5345,95
5346,95
5347,95
5348,95
5349,95
5350,95
5351,95
5352,95
5353,95
5354,95
5355,95
5356,95
5357,95
5358,95
5359,95
5360,95
5361,95
5362,95
5363,95
5364,95
5365,95
5366,95
5367,95
5368,95
5369,95
5370,95
5371,95
5372,95
5373,95
5374,95
5375,95
5376,96
5377,96
5378,96
5379,96
5380,96
5381,96
5382,96
5383,96
5384,96
5385,96
5386,96
5387,96
5388,96
5389,96
5390,96
5391,96
5392,96
5393,96
5394,96
5395,96
5396,96
5397,96
5398,96
5399,96
5400,96
5401,96
5402,96
5403,96
5404,96
5405,96
5406,96
5407,96
5408,96
5409,96
5410,96
5411,96
5412,96
5413,96
5414,96
5415,96
5416,96
5417,96
5418,96
5419,96
5420,96
5421,96
5422,96
5423,96
5424,96
5425,96
5426,96
5427,96
5428,96
5429,96
5430,96
5431,96
5432,97
5433,97
5434,97
5435,97
5436,97
5437,97
5438,97
5439,97
5440,97
5441,97
5442,97
5443,97
5444,97
5445,97
5446,97
5447,97
5448,97
5449,97
5450,97
5451,97
5452,97
5453,97
5454,97
5455,97
5456,97
5457,97
5458,97
5459,97
5460,97
5461,97
5462,97
5463,97
5464,97
5465,97
5466,97
5467,97
5468,97
5469,97
5470,97
5471,97
5472,97
5473,97
5474,97
5475,97
5476,97
5477,97
5478,97
5479,97
5480,97
5481,97
5482,97
5483,97
5484,97
5485,97
5486,97
5487,97
5488,98
5489,98
5490,98
5491,98
5492,98
5493,98
5494,98
5495,98
5496,98
5497,98
5498,98
5499,98
5500,98
5501,98
5502,98
5503,98
5504,98
5505,98
5506,98
5507,98
5508,98
5509,98
5510,98
5511,98
5512,98
5513,98
5514,98
5515,98
5516,98
5517,98
5518,98
5519,98
5520,98
5521,98
5522,98
5523,98
5524,98
5525,98
5526,98
5527,98
5528,98
5529,98
5530,98
5531,98
5532,98
5533,98
5534,98
5535,98
5536,98
5537,98
5538,98
5539,98
5540,98
5541,98
5542,98
5543,98
5544,99
5545,99
5546,99
5547,99
5548,99
5549,99
5550,99
5551,99
5552,99
5553,99
5554,99
5555,99
5556,99
5557,99
5558,99
5559,99
5560,99
5561,99
5562,99
5563,99
5564,99
5565,99
5566,99
5567,99
5568,99
5569,99
5570,99
5571,99
5572,99
5573,99
5574,99
5575,99
5576,99
5577,99
5578,99
5579,99
5580,99
5581,99
5582,99
5583,99
5584,99
5585,99
5586,99
5587,99
5588,99
5589,99
5590,99
5591,99
5592,99
5593,99
5594,99
5595,99
5596,99
5597,99
5598,99
5599,99
5600,100
5601,100
5602,100
5603,100
5604,100
5605,100
5606,100
5607,100
5608,100
5609,100
5610,100
5611,100
5612,100
5613,100
5614,100
5615,100
5616,100
5617,100
5618,100
5619,100
5620,100
5621,100
5622,100
5623,100
5624,100
5625,100
5626,100
5627,100
5628,100
5629,100
5630,100
5631,100
5632,100
5633,100
5634,100
5635,100
5636,100
5637,100
5638,100
5639,100
5640,100
5641,100
5642,100
5643,100
5644,100
5645,100
5646,100
5647,100
5648,100
5649,100
5650,100
5651,100
5652,100
5653,100
5654,100
5655,100
5656,101
5657,101
5658,101
5659,101
5660,101
5661,101
5662,101
5663,101
5664,101
5665,101
5666,101
5667,101
5668,101
5669,101
5670,101
5671,101
5672,101
5673,101
5674,101
5675,101
5676,101
5677,101
5678,101
5679,101
5680,101
5681,101
5682,101
5683,101
5684,101
5685,101
5686,101
5687,101
5688,101
5689,101
5690,101
5691,101
5692,101
5693,101
5694,101
5695,101
5696,101
5697,101
5698,101
5699,101
5700,101
5701,101
5702,101
5703,101
5704,101
5705,101
5706,101
5707,101
5708,101
5709,101
5710,101
5711,101
5712,102
5713,102
5714,102
5715,102
5716,102
5717,102
5718,102
5719,102
5720,102
5721,102
5722,102
5723,102
5724,102
5725,102
5726,102
5727,102
5728,102
5729,102
5730,102
5731,102
5732,102
5733,102
5734,102
5735,102
5736,102
5737,102
5738,102
5739,102
5740,102
5741,102
5742,102
5743,102
5744,102
5745,102
5746,102
5747,102
5748,102
5749,102
5750,102
5751,102
5752,102
5753,102
5754,102
5755,102
5756,102
5757,102
5758,102
5759,102
5760,102
5761,102
5762,102
5763,102
5764,102
5765,102
5766,102
5767,102
5768,103
5769,103
5770,103
5771,103
5772,103
5773,103
5774,103
5775,103
5776,103
5777,103
5778,103
5779,103
5780,103
5781,103
5782,103
5783,103
5784,103
5785,103
5786,103
5787,103
5788,103
5789,103
5790,103
5791,103
5792,103
5793,103
5794,103
5795,103
5796,103
5797,103
5798,103
5799,103
5800,103
5801,103
5802,103
5803,103
5804,103
5805,103
5806,103
5807,103
5808,103
5809,103
5810,103
5811,103
5812,103
5813,103
5814,103
5815,103
5816,103
5817,103
5818,103
5819,103
5820,103
5821,103
5822,103
5823,103
5824,104
5825,104
5826,104
5827,104
5828,104
5829,104
5830,104
5831,104
5832,104
5833,104
5834,104
5835,104
5836,104
5837,104
5838,104
5839,104
5840,104
5841,104
5842,104
5843,104
5844,104
5845,104
5846,104
5847,104
5848,104
5849,104
5850,104
5851,104
5852,104
5853,104
5854,104
5855,104
5856,104
5857,104
5858,104
5859,104
5860,104
5861,104
5862,104
5863,104
5864,104
5865,104
5866,104
5867,104
5868,104
5869,104
5870,104
5871,104
5872,104
5873,104
5874,104
5875,104
5876,104
5877,104
5878,104
5879,104
5880,105
5881,105
5882,105
5883,105
5884,105
5885,105
5886,105
5887,105
5888,105
5889,105
5890,105
5891,105
5892,105
5893,105
5894,105
5895,105
5896,105
5897,105
5898,105
5899,105
5900,105
5901,105
5902,105
5903,105
5904,105
5905,105
5906,105
5907,105
5908,105
5909,105
5910,105
5911,105
5912,105
5913,105
5914,105
5915,105
5916,105
5917,105
5918,105
5919,105
5920,105
5921,105
5922,105
5923,105
5924,105
5925,105
5926,105
5927,105
5928,105
5929,105
5930,105
5931,105
5932,105
5933,105
5934,105
5935,105
5936,106
5937,106
5938,106
5939,106
5940,106
5941,106
5942,106
5943,106
5944,106
5945,106
5946,106
5947,106
5948,106
5949,106
5950,106
5951,106
5952,106
5953,106
5954,106
5955,106
5956,106
5957,106
5958,106
5959,106
5960,106
5961,106
5962,106
5963,106
5964,106
5965,106
5966,106
5967,106
5968,106
5969,106
5970,106
5971,106
5972,106
5973,106
5974,106
5975,106
5976,106
5977,106
5978,106
5979,106
5980,106
5981,106
5982,106
5983,106
5984,106
5985,106
5986,106
5987,106
5988,106
5989,106
5990,106
5991,106
5992,107
5993,107
5994,107
5995,107
5996,107
5997,107
5998,107
5999,107
6000,107
6001,107
6002,107
6003,107
6004,107
6005,107
6006,107
6007,107
6008,107
6009,107
6010,107
6011,107
6012,107
6013,107
6014,107
6015,107
6016,107
6017,107
6018,107
6019,107
6020,107
6021,107
6022,107
6023,107
6024,107
6025,107
6026,107
6027,107
6028,107
6029,107
6030,107
6031,107
6032,107
6033,107
6034,107
6035,107
6036,107
6037,107
6038,107
6039,107
6040,107
6041,107
6042,107
6043,107
6044,107
6045,107
6046,107
6047,107
6048,108
6049,108
6050,108
6051,108
6052,108
6053,108
6054,108
6055,108
6056,108
6057,108
6058,108
6059,108
6060,108
6061,108
6062,108
6063,108
6064,108
6065,108
6066,108
6067,108
6068,108
6069,108
6070,108
6071,108
6072,108
6073,108
6074,108
6075,108
6076,108
6077,108
6078,108
6079,108
6080,108
6081,108
6082,108
6083,108
6084,108
6085,108
6086,108
6087,108
6088,108
6089,108
6090,108
6091,108
6092,108
6093,108
6094,108
6095,108
6096,108
6097,108
6098,108
6099,108
6100,108
6101,108
6102,108
6103,108
6104,109
6105,109
6106,109
6107,109
6108,109
6109,109
6110,109
6111,109
6112,109
6113,109
6114,109
6115,109
6116,109
6117,109
6118,109
6119,109
6120,109
6121,109
6122,109
6123,109
6124,109
6125,109
6126,109
6127,109
6128,109
6129,109
6130,109
6131,109
6132,109
6133,109
6134,109
6135,109
6136,109
6137,109
6138,109
6139,109
6140,109
6141,109
6142,109
6143,109
6144,109
6145,109
6146,109
6147,109
6148,109
6149,109
6150,109
6151,109
6152,109
6153,109
6154,109
6155,109
6156,109
6157,109
6158,109
6159,109
6160,110
6161,110
6162,110
6163,110
6164,110
6165,110
6166,110
6167,110
6168,110
6169,110
6170,110
6171,110
6172,110
6173,110
6174,110
6175,110
6176,110
6177,110
6178,110
6179,110
6180,110
6181,110
6182,110
6183,110
6184,110
6185,110
6186,110
6187,110
6188,110
6189,110
6190,110
6191,110
6192,110
6193,110
6194,110
6195,110
6196,110
6197,110
6198,110
6199,110
6200,110
6201,110
6202,110
6203,110
6204,110
6205,110
6206,110
6207,110
6208,110
6209,110
6210,110
6211,110
6212,110
6213,110
6214,110
6215,110
6216,111
6217,111
6218,111
6219,111
6220,111
6221,111
6222,111
6223,111
6224,111
6225,111
6226,111
6227,111
6228,111
6229,111
6230,111
6231,111
6232,111
6233,111
6234,111
6235,111
6236,111
6237,111
6238,111
6239,111
6240,111
6241,111
6242,111
6243,111
6244,111
6245,111
6246,111
6247,111
6248,111
6249,111
6250,111
6251,111
6252,111
6253,111
6254,111
6255,111
6256,111
6257,111
6258,111
6259,111
6260,111
6261,111
6262,111
6263,111
6264,111
6265,111
6266,111
6267,111
6268,111
6269,111
6270,111
6271,111
6272,112
6273,112
6274,112
6275,112
6276,112
6277,112
6278,112
6279,112
6280,112
6281,112
6282,112
6283,112
6284,112
6285,112
6286,112
6287,112
6288,112
6289,112
6290,112
6291,112
6292,112
6293,112
6294,112
6295,112
6296,112
6297,112
6298,112
6299,112
6300,112
6301,112
6302,112
6303,112
6304,112
6305,112
6306,112
6307,112
6308,112
6309,112
6310,112
6311,112
6312,112
6313,112
6314,112
6315,112
6316,112
6317,112
6318,112
6319,112
6320,112
6321,112
6322,112
6323,112
6324,112
6325,112
6326,112
6327,112
6328,113
6329,113
6330,113
6331,113
6332,113
6333,113
6334,113
6335,113
6336,113
6337,113
6338,113
6339,113
6340,113
6341,113
6342,113
6343,113
6344,113
6345,113
6346,113
6347,113
6348,113
6349,113
6350,113
6351,113
6352,113
6353,113
6354,113
6355,113
6356,113
6357,113
6358,113
6359,113
6360,113
6361,113
6362,113
6363,113
6364,113
6365,113
6366,113
6367,113
6368,113
6369,113
6370,113
6371,113
6372,113
6373,113
6374,113
6375,113
6376,113
6377,113
6378,113
6379,113
6380,113
6381,113
6382,113
6383,113
6384,114
6385,114
6386,114
6387,114
6388,114
6389,114
6390,114
6391,114
6392,114
6393,114
6394,114
6395,114
6396,114
6397,114
6398,114
6399,114
6400,114
6401,114
6402,114
6403,114
6404,114
6405,114
6406,114
6407,114
6408,114
6409,114
6410,114
6411,114
6412,114
6413,114
6414,114
6415,114
6416,114
6417,114
6418,114
6419,114
6420,114
6421,114
6422,114
6423,114
6424,114
6425,114
6426,114
6427,114
6428,114
6429,114
6430,114
6431,114
6432,114
6433,114
6434,114
6435,114
6436,114
6437,114
6438,114
6439,114
6440,115
6441,115
6442,115
6443,115
6444,115
6445,115
6446,115
6447,115
6448,115
6449,115
6450,115
6451,115
6452,115
6453,115
6454,115
6455,115
6456,115
6457,115
6458,115
6459,115
6460,115
6461,115
6462,115
6463,115
6464,115
6465,115
6466,115
6467,115
6468,115
6469,115
6470,115
6471,115
6472,115
6473,115
6474,115
6475,115
6476,115
6477,115
6478,115
6479,115
6480,115
6481,115
6482,115
6483,115
6484,115
6485,115
6486,115
6487,115
6488,115
6489,115
6490,115
6491,115
6492,115
6493,115
6494,115
6495,115
6496,116
6497,116
6498,116
6499,116
6500,116
6501,116
6502,116
6503,116
6504,116
6505,116
6506,116
6507,116
6508,116
6509,116
6510,116
6511,116
6512,116
6513,116
6514,116
6515,116
6516,116
6517,116
6518,116
6519,116
6520,116
6521,116
6522,116
6523,116
6524,116
6525,116
6526,116
6527,116
6528,116
6529,116
6530,116
6531,116
6532,116
6533,116
6534,116
6535,116
6536,116
6537,116
6538,116
6539,116
6540,116
6541,116
6542,116
6543,116
6544,116
6545,116
6546,116
6547,116
6548,116
6549,116
6550,116
6551,116
6552,117
6553,117
6554,117
6555,117
6556,117
6557,117
6558,117
6559,117
6560,117
6561,117
6562,117
6563,117
6564,117
6565,117
6566,117
6567,117
6568,117
6569,117
6570,117
6571,117
6572,117
6573,117
6574,117
6575,117
6576,117
6577,117
6578,117
6579,117
6580,117
6581,117
6582,117
6583,117
6584,117
6585,117
6586,117
6587,117
6588,117
6589,117
6590,117
6591,117
6592,117
6593,117
6594,117
6595,117
6596,117
6597,117
6598,117
6599,117
6600,117
6601,117
6602,117
6603,117
6604,117
6605,117
6606,117
6607,117
6608,118
6609,118
6610,118
6611,118
6612,118
6613,118
6614,118
6615,118
6616,118
6617,118
6618,118
6619,118
6620,118
6621,118
6622,118
6623,118
6624,118
6625,118
6626,118
6627,118
6628,118
6629,118
6630,118
6631,118
6632,118
6633,118
6634,118
6635,118
6636,118
6637,118
6638,118
6639,118
6640,118
6641,118
6642,118
6643,118
6644,118
6645,118
6646,118
6647,118
6648,118
6649,118
6650,118
6651,118
6652,118
6653,118
6654,118
6655,118
6656,118
6657,118
6658,118
6659,118
6660,118
6661,118
6662,118
6663,118
6664,119
6665,119
6666,119
6667,119
6668,119
6669,119
6670,119
6671,119
6672,119
6673,119
6674,119
6675,119
6676,119
6677,119
6678,119
6679,119
6680,119
6681,119
6682,119
6683,119
6684,119
6685,119
6686,119
6687,119
6688,119
6689,119
6690,119
6691,119
6692,119
6693,119
6694,119
6695,119
6696,119
6697,119
6698,119
6699,119
6700,119
6701,119
6702,119
6703,119
6704,119
6705,119
6706,119
6707,119
6708,119
6709,119
6710,119
6711,119
6712,119
6713,119
6714,119
6715,119
6716,119
6717,119
6718,119
6719,119
