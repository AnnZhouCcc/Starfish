0,0
1,0
2,0
3,0
4,0
5,0
6,0
7,0
8,0
9,0
10,0
11,0
12,0
13,0
14,0
15,0
16,0
17,0
18,0
19,0
20,0
21,0
22,0
23,0
24,0
25,0
26,0
27,0
28,1
29,1
30,1
31,1
32,1
33,1
34,1
35,1
36,1
37,1
38,1
39,1
40,1
41,1
42,1
43,1
44,1
45,1
46,1
47,1
48,1
49,1
50,1
51,1
52,1
53,1
54,1
55,1
56,2
57,2
58,2
59,2
60,2
61,2
62,2
63,2
64,2
65,2
66,2
67,2
68,2
69,2
70,2
71,2
72,2
73,2
74,2
75,2
76,2
77,2
78,2
79,2
80,2
81,2
82,2
83,2
84,3
85,3
86,3
87,3
88,3
89,3
90,3
91,3
92,3
93,3
94,3
95,3
96,3
97,3
98,3
99,3
100,3
101,3
102,3
103,3
104,3
105,3
106,3
107,3
108,3
109,3
110,3
111,3
112,4
113,4
114,4
115,4
116,4
117,4
118,4
119,4
120,4
121,4
122,4
123,4
124,4
125,4
126,4
127,4
128,4
129,4
130,4
131,4
132,4
133,4
134,4
135,4
136,4
137,4
138,4
139,4
140,5
141,5
142,5
143,5
144,5
145,5
146,5
147,5
148,5
149,5
150,5
151,5
152,5
153,5
154,5
155,5
156,5
157,5
158,5
159,5
160,5
161,5
162,5
163,5
164,5
165,5
166,5
167,5
168,6
169,6
170,6
171,6
172,6
173,6
174,6
175,6
176,6
177,6
178,6
179,6
180,6
181,6
182,6
183,6
184,6
185,6
186,6
187,6
188,6
189,6
190,6
191,6
192,6
193,6
194,6
195,6
196,7
197,7
198,7
199,7
200,7
201,7
202,7
203,7
204,7
205,7
206,7
207,7
208,7
209,7
210,7
211,7
212,7
213,7
214,7
215,7
216,7
217,7
218,7
219,7
220,7
221,7
222,7
223,7
224,8
225,8
226,8
227,8
228,8
229,8
230,8
231,8
232,8
233,8
234,8
235,8
236,8
237,8
238,8
239,8
240,8
241,8
242,8
243,8
244,8
245,8
246,8
247,8
248,8
249,8
250,8
251,8
252,9
253,9
254,9
255,9
256,9
257,9
258,9
259,9
260,9
261,9
262,9
263,9
264,9
265,9
266,9
267,9
268,9
269,9
270,9
271,9
272,9
273,9
274,9
275,9
276,9
277,9
278,9
279,9
280,10
281,10
282,10
283,10
284,10
285,10
286,10
287,10
288,10
289,10
290,10
291,10
292,10
293,10
294,10
295,10
296,10
297,10
298,10
299,10
300,10
301,10
302,10
303,10
304,10
305,10
306,10
307,10
308,11
309,11
310,11
311,11
312,11
313,11
314,11
315,11
316,11
317,11
318,11
319,11
320,11
321,11
322,11
323,11
324,11
325,11
326,11
327,11
328,11
329,11
330,11
331,11
332,11
333,11
334,11
335,11
336,12
337,12
338,12
339,12
340,12
341,12
342,12
343,12
344,12
345,12
346,12
347,12
348,12
349,12
350,12
351,12
352,12
353,12
354,12
355,12
356,12
357,12
358,12
359,12
360,12
361,12
362,12
363,12
364,13
365,13
366,13
367,13
368,13
369,13
370,13
371,13
372,13
373,13
374,13
375,13
376,13
377,13
378,13
379,13
380,13
381,13
382,13
383,13
384,13
385,13
386,13
387,13
388,13
389,13
390,13
391,13
392,14
393,14
394,14
395,14
396,14
397,14
398,14
399,14
400,14
401,14
402,14
403,14
404,14
405,14
406,14
407,14
408,14
409,14
410,14
411,14
412,14
413,14
414,14
415,14
416,14
417,14
418,14
419,14
420,15
421,15
422,15
423,15
424,15
425,15
426,15
427,15
428,15
429,15
430,15
431,15
432,15
433,15
434,15
435,15
436,15
437,15
438,15
439,15
440,15
441,15
442,15
443,15
444,15
445,15
446,15
447,15
448,16
449,16
450,16
451,16
452,16
453,16
454,16
455,16
456,16
457,16
458,16
459,16
460,16
461,16
462,16
463,16
464,16
465,16
466,16
467,16
468,16
469,16
470,16
471,16
472,16
473,16
474,16
475,16
476,17
477,17
478,17
479,17
480,17
481,17
482,17
483,17
484,17
485,17
486,17
487,17
488,17
489,17
490,17
491,17
492,17
493,17
494,17
495,17
496,17
497,17
498,17
499,17
500,17
501,17
502,17
503,17
504,18
505,18
506,18
507,18
508,18
509,18
510,18
511,18
512,18
513,18
514,18
515,18
516,18
517,18
518,18
519,18
520,18
521,18
522,18
523,18
524,18
525,18
526,18
527,18
528,18
529,18
530,18
531,18
532,19
533,19
534,19
535,19
536,19
537,19
538,19
539,19
540,19
541,19
542,19
543,19
544,19
545,19
546,19
547,19
548,19
549,19
550,19
551,19
552,19
553,19
554,19
555,19
556,19
557,19
558,19
559,19
560,20
561,20
562,20
563,20
564,20
565,20
566,20
567,20
568,20
569,20
570,20
571,20
572,20
573,20
574,20
575,20
576,20
577,20
578,20
579,20
580,20
581,20
582,20
583,20
584,20
585,20
586,20
587,20
588,21
589,21
590,21
591,21
592,21
593,21
594,21
595,21
596,21
597,21
598,21
599,21
600,21
601,21
602,21
603,21
604,21
605,21
606,21
607,21
608,21
609,21
610,21
611,21
612,21
613,21
614,21
615,21
616,22
617,22
618,22
619,22
620,22
621,22
622,22
623,22
624,22
625,22
626,22
627,22
628,22
629,22
630,22
631,22
632,22
633,22
634,22
635,22
636,22
637,22
638,22
639,22
640,22
641,22
642,22
643,22
644,23
645,23
646,23
647,23
648,23
649,23
650,23
651,23
652,23
653,23
654,23
655,23
656,23
657,23
658,23
659,23
660,23
661,23
662,23
663,23
664,23
665,23
666,23
667,23
668,23
669,23
670,23
671,23
672,24
673,24
674,24
675,24
676,24
677,24
678,24
679,24
680,24
681,24
682,24
683,24
684,24
685,24
686,24
687,24
688,24
689,24
690,24
691,24
692,24
693,24
694,24
695,24
696,24
697,24
698,24
699,24
700,25
701,25
702,25
703,25
704,25
705,25
706,25
707,25
708,25
709,25
710,25
711,25
712,25
713,25
714,25
715,25
716,25
717,25
718,25
719,25
720,25
721,25
722,25
723,25
724,25
725,25
726,25
727,25
728,26
729,26
730,26
731,26
732,26
733,26
734,26
735,26
736,26
737,26
738,26
739,26
740,26
741,26
742,26
743,26
744,26
745,26
746,26
747,26
748,26
749,26
750,26
751,26
752,26
753,26
754,26
755,26
756,27
757,27
758,27
759,27
760,27
761,27
762,27
763,27
764,27
765,27
766,27
767,27
768,27
769,27
770,27
771,27
772,27
773,27
774,27
775,27
776,27
777,27
778,27
779,27
780,27
781,27
782,27
783,27
784,28
785,28
786,28
787,28
788,28
789,28
790,28
791,28
792,28
793,28
794,28
795,28
796,28
797,28
798,28
799,28
800,28
801,28
802,28
803,28
804,28
805,28
806,28
807,28
808,28
809,28
810,28
811,28
812,29
813,29
814,29
815,29
816,29
817,29
818,29
819,29
820,29
821,29
822,29
823,29
824,29
825,29
826,29
827,29
828,29
829,29
830,29
831,29
832,29
833,29
834,29
835,29
836,29
837,29
838,29
839,29
840,30
841,30
842,30
843,30
844,30
845,30
846,30
847,30
848,30
849,30
850,30
851,30
852,30
853,30
854,30
855,30
856,30
857,30
858,30
859,30
860,30
861,30
862,30
863,30
864,30
865,30
866,30
867,30
868,31
869,31
870,31
871,31
872,31
873,31
874,31
875,31
876,31
877,31
878,31
879,31
880,31
881,31
882,31
883,31
884,31
885,31
886,31
887,31
888,31
889,31
890,31
891,31
892,31
893,31
894,31
895,31
896,32
897,32
898,32
899,32
900,32
901,32
902,32
903,32
904,32
905,32
906,32
907,32
908,32
909,32
910,32
911,32
912,32
913,32
914,32
915,32
916,32
917,32
918,32
919,32
920,32
921,32
922,32
923,32
924,33
925,33
926,33
927,33
928,33
929,33
930,33
931,33
932,33
933,33
934,33
935,33
936,33
937,33
938,33
939,33
940,33
941,33
942,33
943,33
944,33
945,33
946,33
947,33
948,33
949,33
950,33
951,33
952,34
953,34
954,34
955,34
956,34
957,34
958,34
959,34
960,34
961,34
962,34
963,34
964,34
965,34
966,34
967,34
968,34
969,34
970,34
971,34
972,34
973,34
974,34
975,34
976,34
977,34
978,34
979,34
980,35
981,35
982,35
983,35
984,35
985,35
986,35
987,35
988,35
989,35
990,35
991,35
992,35
993,35
994,35
995,35
996,35
997,35
998,35
999,35
1000,35
1001,35
1002,35
1003,35
1004,35
1005,35
1006,35
1007,35
1008,36
1009,36
1010,36
1011,36
1012,36
1013,36
1014,36
1015,36
1016,36
1017,36
1018,36
1019,36
1020,36
1021,36
1022,36
1023,36
1024,36
1025,36
1026,36
1027,36
1028,36
1029,36
1030,36
1031,36
1032,36
1033,36
1034,36
1035,36
1036,37
1037,37
1038,37
1039,37
1040,37
1041,37
1042,37
1043,37
1044,37
1045,37
1046,37
1047,37
1048,37
1049,37
1050,37
1051,37
1052,37
1053,37
1054,37
1055,37
1056,37
1057,37
1058,37
1059,37
1060,37
1061,37
1062,37
1063,37
1064,38
1065,38
1066,38
1067,38
1068,38
1069,38
1070,38
1071,38
1072,38
1073,38
1074,38
1075,38
1076,38
1077,38
1078,38
1079,38
1080,38
1081,38
1082,38
1083,38
1084,38
1085,38
1086,38
1087,38
1088,38
1089,38
1090,38
1091,38
1092,39
1093,39
1094,39
1095,39
1096,39
1097,39
1098,39
1099,39
1100,39
1101,39
1102,39
1103,39
1104,39
1105,39
1106,39
1107,39
1108,39
1109,39
1110,39
1111,39
1112,39
1113,39
1114,39
1115,39
1116,39
1117,39
1118,39
1119,39
1120,40
1121,40
1122,40
1123,40
1124,40
1125,40
1126,40
1127,40
1128,40
1129,40
1130,40
1131,40
1132,40
1133,40
1134,40
1135,40
1136,40
1137,40
1138,40
1139,40
1140,40
1141,40
1142,40
1143,40
1144,40
1145,40
1146,40
1147,40
1148,41
1149,41
1150,41
1151,41
1152,41
1153,41
1154,41
1155,41
1156,41
1157,41
1158,41
1159,41
1160,41
1161,41
1162,41
1163,41
1164,41
1165,41
1166,41
1167,41
1168,41
1169,41
1170,41
1171,41
1172,41
1173,41
1174,41
1175,41
1176,42
1177,42
1178,42
1179,42
1180,42
1181,42
1182,42
1183,42
1184,42
1185,42
1186,42
1187,42
1188,42
1189,42
1190,42
1191,42
1192,42
1193,42
1194,42
1195,42
1196,42
1197,42
1198,42
1199,42
1200,42
1201,42
1202,42
1203,42
1204,43
1205,43
1206,43
1207,43
1208,43
1209,43
1210,43
1211,43
1212,43
1213,43
1214,43
1215,43
1216,43
1217,43
1218,43
1219,43
1220,43
1221,43
1222,43
1223,43
1224,43
1225,43
1226,43
1227,43
1228,43
1229,43
1230,43
1231,43
1232,44
1233,44
1234,44
1235,44
1236,44
1237,44
1238,44
1239,44
1240,44
1241,44
1242,44
1243,44
1244,44
1245,44
1246,44
1247,44
1248,44
1249,44
1250,44
1251,44
1252,44
1253,44
1254,44
1255,44
1256,44
1257,44
1258,44
1259,44
1260,45
1261,45
1262,45
1263,45
1264,45
1265,45
1266,45
1267,45
1268,45
1269,45
1270,45
1271,45
1272,45
1273,45
1274,45
1275,45
1276,45
1277,45
1278,45
1279,45
1280,45
1281,45
1282,45
1283,45
1284,45
1285,45
1286,45
1287,45
1288,46
1289,46
1290,46
1291,46
1292,46
1293,46
1294,46
1295,46
1296,46
1297,46
1298,46
1299,46
1300,46
1301,46
1302,46
1303,46
1304,46
1305,46
1306,46
1307,46
1308,46
1309,46
1310,46
1311,46
1312,46
1313,46
1314,46
1315,46
1316,47
1317,47
1318,47
1319,47
1320,47
1321,47
1322,47
1323,47
1324,47
1325,47
1326,47
1327,47
1328,47
1329,47
1330,47
1331,47
1332,47
1333,47
1334,47
1335,47
1336,47
1337,47
1338,47
1339,47
1340,47
1341,47
1342,47
1343,47
1344,48
1345,48
1346,48
1347,48
1348,48
1349,48
1350,48
1351,48
1352,48
1353,48
1354,48
1355,48
1356,48
1357,48
1358,48
1359,48
1360,48
1361,48
1362,48
1363,48
1364,48
1365,48
1366,48
1367,48
1368,48
1369,48
1370,48
1371,48
1372,49
1373,49
1374,49
1375,49
1376,49
1377,49
1378,49
1379,49
1380,49
1381,49
1382,49
1383,49
1384,49
1385,49
1386,49
1387,49
1388,49
1389,49
1390,49
1391,49
1392,49
1393,49
1394,49
1395,49
1396,49
1397,49
1398,49
1399,49
1400,50
1401,50
1402,50
1403,50
1404,50
1405,50
1406,50
1407,50
1408,50
1409,50
1410,50
1411,50
1412,50
1413,50
1414,50
1415,50
1416,50
1417,50
1418,50
1419,50
1420,50
1421,50
1422,50
1423,50
1424,50
1425,50
1426,50
1427,50
1428,51
1429,51
1430,51
1431,51
1432,51
1433,51
1434,51
1435,51
1436,51
1437,51
1438,51
1439,51
1440,51
1441,51
1442,51
1443,51
1444,51
1445,51
1446,51
1447,51
1448,51
1449,51
1450,51
1451,51
1452,51
1453,51
1454,51
1455,51
1456,52
1457,52
1458,52
1459,52
1460,52
1461,52
1462,52
1463,52
1464,52
1465,52
1466,52
1467,52
1468,52
1469,52
1470,52
1471,52
1472,52
1473,52
1474,52
1475,52
1476,52
1477,52
1478,52
1479,52
1480,52
1481,52
1482,52
1483,52
1484,53
1485,53
1486,53
1487,53
1488,53
1489,53
1490,53
1491,53
1492,53
1493,53
1494,53
1495,53
1496,53
1497,53
1498,53
1499,53
1500,53
1501,53
1502,53
1503,53
1504,53
1505,53
1506,53
1507,53
1508,53
1509,53
1510,53
1511,53
1512,54
1513,54
1514,54
1515,54
1516,54
1517,54
1518,54
1519,54
1520,54
1521,54
1522,54
1523,54
1524,54
1525,54
1526,54
1527,54
1528,54
1529,54
1530,54
1531,54
1532,54
1533,54
1534,54
1535,54
1536,54
1537,54
1538,54
1539,54
1540,55
1541,55
1542,55
1543,55
1544,55
1545,55
1546,55
1547,55
1548,55
1549,55
1550,55
1551,55
1552,55
1553,55
1554,55
1555,55
1556,55
1557,55
1558,55
1559,55
1560,55
1561,55
1562,55
1563,55
1564,55
1565,55
1566,55
1567,55
1568,56
1569,56
1570,56
1571,56
1572,56
1573,56
1574,56
1575,56
1576,56
1577,56
1578,56
1579,56
1580,56
1581,56
1582,56
1583,56
1584,56
1585,56
1586,56
1587,56
1588,56
1589,56
1590,56
1591,56
1592,56
1593,56
1594,56
1595,56
1596,57
1597,57
1598,57
1599,57
1600,57
1601,57
1602,57
1603,57
1604,57
1605,57
1606,57
1607,57
1608,57
1609,57
1610,57
1611,57
1612,57
1613,57
1614,57
1615,57
1616,57
1617,57
1618,57
1619,57
1620,57
1621,57
1622,57
1623,57
1624,58
1625,58
1626,58
1627,58
1628,58
1629,58
1630,58
1631,58
1632,58
1633,58
1634,58
1635,58
1636,58
1637,58
1638,58
1639,58
1640,58
1641,58
1642,58
1643,58
1644,58
1645,58
1646,58
1647,58
1648,58
1649,58
1650,58
1651,58
1652,59
1653,59
1654,59
1655,59
1656,59
1657,59
1658,59
1659,59
1660,59
1661,59
1662,59
1663,59
1664,59
1665,59
1666,59
1667,59
1668,59
1669,59
1670,59
1671,59
1672,59
1673,59
1674,59
1675,59
1676,59
1677,59
1678,59
1679,59
