0,0
1,0
2,0
3,0
4,0
5,0
6,0
7,0
8,0
9,0
10,0
11,0
12,0
13,0
14,0
15,0
16,0
17,0
18,0
19,0
20,0
21,0
22,0
23,0
24,0
25,0
26,0
27,0
28,0
29,0
30,0
31,0
32,0
33,0
34,0
35,0
36,0
37,0
38,0
39,0
40,1
41,1
42,1
43,1
44,1
45,1
46,1
47,1
48,1
49,1
50,1
51,1
52,1
53,1
54,1
55,1
56,1
57,1
58,1
59,1
60,1
61,1
62,1
63,1
64,1
65,1
66,1
67,1
68,1
69,1
70,1
71,1
72,1
73,1
74,1
75,1
76,1
77,1
78,1
79,1
80,2
81,2
82,2
83,2
84,2
85,2
86,2
87,2
88,2
89,2
90,2
91,2
92,2
93,2
94,2
95,2
96,2
97,2
98,2
99,2
100,2
101,2
102,2
103,2
104,2
105,2
106,2
107,2
108,2
109,2
110,2
111,2
112,2
113,2
114,2
115,2
116,2
117,2
118,2
119,2
120,3
121,3
122,3
123,3
124,3
125,3
126,3
127,3
128,3
129,3
130,3
131,3
132,3
133,3
134,3
135,3
136,3
137,3
138,3
139,3
140,3
141,3
142,3
143,3
144,3
145,3
146,3
147,3
148,3
149,3
150,3
151,3
152,3
153,3
154,3
155,3
156,3
157,3
158,3
159,3
160,4
161,4
162,4
163,4
164,4
165,4
166,4
167,4
168,4
169,4
170,4
171,4
172,4
173,4
174,4
175,4
176,4
177,4
178,4
179,4
180,4
181,4
182,4
183,4
184,4
185,4
186,4
187,4
188,4
189,4
190,4
191,4
192,4
193,4
194,4
195,4
196,4
197,4
198,4
199,4
200,5
201,5
202,5
203,5
204,5
205,5
206,5
207,5
208,5
209,5
210,5
211,5
212,5
213,5
214,5
215,5
216,5
217,5
218,5
219,5
220,5
221,5
222,5
223,5
224,5
225,5
226,5
227,5
228,5
229,5
230,5
231,5
232,5
233,5
234,5
235,5
236,5
237,5
238,5
239,5
240,6
241,6
242,6
243,6
244,6
245,6
246,6
247,6
248,6
249,6
250,6
251,6
252,6
253,6
254,6
255,6
256,6
257,6
258,6
259,6
260,6
261,6
262,6
263,6
264,6
265,6
266,6
267,6
268,6
269,6
270,6
271,6
272,6
273,6
274,6
275,6
276,6
277,6
278,6
279,6
280,7
281,7
282,7
283,7
284,7
285,7
286,7
287,7
288,7
289,7
290,7
291,7
292,7
293,7
294,7
295,7
296,7
297,7
298,7
299,7
300,7
301,7
302,7
303,7
304,7
305,7
306,7
307,7
308,7
309,7
310,7
311,7
312,7
313,7
314,7
315,7
316,7
317,7
318,7
319,7
320,8
321,8
322,8
323,8
324,8
325,8
326,8
327,8
328,8
329,8
330,8
331,8
332,8
333,8
334,8
335,8
336,8
337,8
338,8
339,8
340,8
341,8
342,8
343,8
344,8
345,8
346,8
347,8
348,8
349,8
350,8
351,8
352,8
353,8
354,8
355,8
356,8
357,8
358,8
359,8
360,9
361,9
362,9
363,9
364,9
365,9
366,9
367,9
368,9
369,9
370,9
371,9
372,9
373,9
374,9
375,9
376,9
377,9
378,9
379,9
380,9
381,9
382,9
383,9
384,9
385,9
386,9
387,9
388,9
389,9
390,9
391,9
392,9
393,9
394,9
395,9
396,9
397,9
398,9
399,9
400,10
401,10
402,10
403,10
404,10
405,10
406,10
407,10
408,10
409,10
410,10
411,10
412,10
413,10
414,10
415,10
416,10
417,10
418,10
419,10
420,10
421,10
422,10
423,10
424,10
425,10
426,10
427,10
428,10
429,10
430,10
431,10
432,10
433,10
434,10
435,10
436,10
437,10
438,10
439,10
440,11
441,11
442,11
443,11
444,11
445,11
446,11
447,11
448,11
449,11
450,11
451,11
452,11
453,11
454,11
455,11
456,11
457,11
458,11
459,11
460,11
461,11
462,11
463,11
464,11
465,11
466,11
467,11
468,11
469,11
470,11
471,11
472,11
473,11
474,11
475,11
476,11
477,11
478,11
479,11
480,12
481,12
482,12
483,12
484,12
485,12
486,12
487,12
488,12
489,12
490,12
491,12
492,12
493,12
494,12
495,12
496,12
497,12
498,12
499,12
500,12
501,12
502,12
503,12
504,12
505,12
506,12
507,12
508,12
509,12
510,12
511,12
512,12
513,12
514,12
515,12
516,12
517,12
518,12
519,12
520,13
521,13
522,13
523,13
524,13
525,13
526,13
527,13
528,13
529,13
530,13
531,13
532,13
533,13
534,13
535,13
536,13
537,13
538,13
539,13
540,13
541,13
542,13
543,13
544,13
545,13
546,13
547,13
548,13
549,13
550,13
551,13
552,13
553,13
554,13
555,13
556,13
557,13
558,13
559,13
560,14
561,14
562,14
563,14
564,14
565,14
566,14
567,14
568,14
569,14
570,14
571,14
572,14
573,14
574,14
575,14
576,14
577,14
578,14
579,14
580,14
581,14
582,14
583,14
584,14
585,14
586,14
587,14
588,14
589,14
590,14
591,14
592,14
593,14
594,14
595,14
596,14
597,14
598,14
599,14
600,15
601,15
602,15
603,15
604,15
605,15
606,15
607,15
608,15
609,15
610,15
611,15
612,15
613,15
614,15
615,15
616,15
617,15
618,15
619,15
620,15
621,15
622,15
623,15
624,15
625,15
626,15
627,15
628,15
629,15
630,15
631,15
632,15
633,15
634,15
635,15
636,15
637,15
638,15
639,15
640,16
641,16
642,16
643,16
644,16
645,16
646,16
647,16
648,16
649,16
650,16
651,16
652,16
653,16
654,16
655,16
656,16
657,16
658,16
659,16
660,16
661,16
662,16
663,16
664,16
665,16
666,16
667,16
668,16
669,16
670,16
671,16
672,16
673,16
674,16
675,16
676,16
677,16
678,16
679,16
680,17
681,17
682,17
683,17
684,17
685,17
686,17
687,17
688,17
689,17
690,17
691,17
692,17
693,17
694,17
695,17
696,17
697,17
698,17
699,17
700,17
701,17
702,17
703,17
704,17
705,17
706,17
707,17
708,17
709,17
710,17
711,17
712,17
713,17
714,17
715,17
716,17
717,17
718,17
719,17
720,18
721,18
722,18
723,18
724,18
725,18
726,18
727,18
728,18
729,18
730,18
731,18
732,18
733,18
734,18
735,18
736,18
737,18
738,18
739,18
740,18
741,18
742,18
743,18
744,18
745,18
746,18
747,18
748,18
749,18
750,18
751,18
752,18
753,18
754,18
755,18
756,18
757,18
758,18
759,18
760,19
761,19
762,19
763,19
764,19
765,19
766,19
767,19
768,19
769,19
770,19
771,19
772,19
773,19
774,19
775,19
776,19
777,19
778,19
779,19
780,19
781,19
782,19
783,19
784,19
785,19
786,19
787,19
788,19
789,19
790,19
791,19
792,19
793,19
794,19
795,19
796,19
797,19
798,19
799,19
800,20
801,20
802,20
803,20
804,20
805,20
806,20
807,20
808,20
809,20
810,20
811,20
812,20
813,20
814,20
815,20
816,20
817,20
818,20
819,20
820,20
821,20
822,20
823,20
824,20
825,20
826,20
827,20
828,20
829,20
830,20
831,20
832,20
833,20
834,20
835,20
836,20
837,20
838,20
839,20
840,21
841,21
842,21
843,21
844,21
845,21
846,21
847,21
848,21
849,21
850,21
851,21
852,21
853,21
854,21
855,21
856,21
857,21
858,21
859,21
860,21
861,21
862,21
863,21
864,21
865,21
866,21
867,21
868,21
869,21
870,21
871,21
872,21
873,21
874,21
875,21
876,21
877,21
878,21
879,21
880,22
881,22
882,22
883,22
884,22
885,22
886,22
887,22
888,22
889,22
890,22
891,22
892,22
893,22
894,22
895,22
896,22
897,22
898,22
899,22
900,22
901,22
902,22
903,22
904,22
905,22
906,22
907,22
908,22
909,22
910,22
911,22
912,22
913,22
914,22
915,22
916,22
917,22
918,22
919,22
920,23
921,23
922,23
923,23
924,23
925,23
926,23
927,23
928,23
929,23
930,23
931,23
932,23
933,23
934,23
935,23
936,23
937,23
938,23
939,23
940,23
941,23
942,23
943,23
944,23
945,23
946,23
947,23
948,23
949,23
950,23
951,23
952,23
953,23
954,23
955,23
956,23
957,23
958,23
959,23
960,24
961,24
962,24
963,24
964,24
965,24
966,24
967,24
968,24
969,24
970,24
971,24
972,24
973,24
974,24
975,24
976,24
977,24
978,24
979,24
980,24
981,24
982,24
983,24
984,24
985,24
986,24
987,24
988,24
989,24
990,24
991,24
992,24
993,24
994,24
995,24
996,24
997,24
998,24
999,24
1000,25
1001,25
1002,25
1003,25
1004,25
1005,25
1006,25
1007,25
1008,25
1009,25
1010,25
1011,25
1012,25
1013,25
1014,25
1015,25
1016,25
1017,25
1018,25
1019,25
1020,25
1021,25
1022,25
1023,25
1024,25
1025,25
1026,25
1027,25
1028,25
1029,25
1030,25
1031,25
1032,25
1033,25
1034,25
1035,25
1036,25
1037,25
1038,25
1039,25
1040,26
1041,26
1042,26
1043,26
1044,26
1045,26
1046,26
1047,26
1048,26
1049,26
1050,26
1051,26
1052,26
1053,26
1054,26
1055,26
1056,26
1057,26
1058,26
1059,26
1060,26
1061,26
1062,26
1063,26
1064,26
1065,26
1066,26
1067,26
1068,26
1069,26
1070,26
1071,26
1072,26
1073,26
1074,26
1075,26
1076,26
1077,26
1078,26
1079,26
1080,27
1081,27
1082,27
1083,27
1084,27
1085,27
1086,27
1087,27
1088,27
1089,27
1090,27
1091,27
1092,27
1093,27
1094,27
1095,27
1096,27
1097,27
1098,27
1099,27
1100,27
1101,27
1102,27
1103,27
1104,27
1105,27
1106,27
1107,27
1108,27
1109,27
1110,27
1111,27
1112,27
1113,27
1114,27
1115,27
1116,27
1117,27
1118,27
1119,27
1120,28
1121,28
1122,28
1123,28
1124,28
1125,28
1126,28
1127,28
1128,28
1129,28
1130,28
1131,28
1132,28
1133,28
1134,28
1135,28
1136,28
1137,28
1138,28
1139,28
1140,28
1141,28
1142,28
1143,28
1144,28
1145,28
1146,28
1147,28
1148,28
1149,28
1150,28
1151,28
1152,28
1153,28
1154,28
1155,28
1156,28
1157,28
1158,28
1159,28
1160,29
1161,29
1162,29
1163,29
1164,29
1165,29
1166,29
1167,29
1168,29
1169,29
1170,29
1171,29
1172,29
1173,29
1174,29
1175,29
1176,29
1177,29
1178,29
1179,29
1180,29
1181,29
1182,29
1183,29
1184,29
1185,29
1186,29
1187,29
1188,29
1189,29
1190,29
1191,29
1192,29
1193,29
1194,29
1195,29
1196,29
1197,29
1198,29
1199,29
1200,30
1201,30
1202,30
1203,30
1204,30
1205,30
1206,30
1207,30
1208,30
1209,30
1210,30
1211,30
1212,30
1213,30
1214,30
1215,30
1216,30
1217,30
1218,30
1219,30
1220,30
1221,30
1222,30
1223,30
1224,30
1225,30
1226,30
1227,30
1228,30
1229,30
1230,30
1231,30
1232,30
1233,30
1234,30
1235,30
1236,30
1237,30
1238,30
1239,30
1240,31
1241,31
1242,31
1243,31
1244,31
1245,31
1246,31
1247,31
1248,31
1249,31
1250,31
1251,31
1252,31
1253,31
1254,31
1255,31
1256,31
1257,31
1258,31
1259,31
1260,31
1261,31
1262,31
1263,31
1264,31
1265,31
1266,31
1267,31
1268,31
1269,31
1270,31
1271,31
1272,31
1273,31
1274,31
1275,31
1276,31
1277,31
1278,31
1279,31
1280,32
1281,32
1282,32
1283,32
1284,32
1285,32
1286,32
1287,32
1288,32
1289,32
1290,32
1291,32
1292,32
1293,32
1294,32
1295,32
1296,32
1297,32
1298,32
1299,32
1300,32
1301,32
1302,32
1303,32
1304,32
1305,32
1306,32
1307,32
1308,32
1309,32
1310,32
1311,32
1312,32
1313,32
1314,32
1315,32
1316,32
1317,32
1318,32
1319,32
1320,33
1321,33
1322,33
1323,33
1324,33
1325,33
1326,33
1327,33
1328,33
1329,33
1330,33
1331,33
1332,33
1333,33
1334,33
1335,33
1336,33
1337,33
1338,33
1339,33
1340,33
1341,33
1342,33
1343,33
1344,33
1345,33
1346,33
1347,33
1348,33
1349,33
1350,33
1351,33
1352,33
1353,33
1354,33
1355,33
1356,33
1357,33
1358,33
1359,33
1360,34
1361,34
1362,34
1363,34
1364,34
1365,34
1366,34
1367,34
1368,34
1369,34
1370,34
1371,34
1372,34
1373,34
1374,34
1375,34
1376,34
1377,34
1378,34
1379,34
1380,34
1381,34
1382,34
1383,34
1384,34
1385,34
1386,34
1387,34
1388,34
1389,34
1390,34
1391,34
1392,34
1393,34
1394,34
1395,34
1396,34
1397,34
1398,34
1399,34
1400,35
1401,35
1402,35
1403,35
1404,35
1405,35
1406,35
1407,35
1408,35
1409,35
1410,35
1411,35
1412,35
1413,35
1414,35
1415,35
1416,35
1417,35
1418,35
1419,35
1420,35
1421,35
1422,35
1423,35
1424,35
1425,35
1426,35
1427,35
1428,35
1429,35
1430,35
1431,35
1432,35
1433,35
1434,35
1435,35
1436,35
1437,35
1438,35
1439,35
1440,36
1441,36
1442,36
1443,36
1444,36
1445,36
1446,36
1447,36
1448,36
1449,36
1450,36
1451,36
1452,36
1453,36
1454,36
1455,36
1456,36
1457,36
1458,36
1459,36
1460,36
1461,36
1462,36
1463,36
1464,36
1465,36
1466,36
1467,36
1468,36
1469,36
1470,36
1471,36
1472,36
1473,36
1474,36
1475,36
1476,36
1477,36
1478,36
1479,36
1480,37
1481,37
1482,37
1483,37
1484,37
1485,37
1486,37
1487,37
1488,37
1489,37
1490,37
1491,37
1492,37
1493,37
1494,37
1495,37
1496,37
1497,37
1498,37
1499,37
1500,37
1501,37
1502,37
1503,37
1504,37
1505,37
1506,37
1507,37
1508,37
1509,37
1510,37
1511,37
1512,37
1513,37
1514,37
1515,37
1516,37
1517,37
1518,37
1519,37
1520,38
1521,38
1522,38
1523,38
1524,38
1525,38
1526,38
1527,38
1528,38
1529,38
1530,38
1531,38
1532,38
1533,38
1534,38
1535,38
1536,38
1537,38
1538,38
1539,38
1540,38
1541,38
1542,38
1543,38
1544,38
1545,38
1546,38
1547,38
1548,38
1549,38
1550,38
1551,38
1552,38
1553,38
1554,38
1555,38
1556,38
1557,38
1558,38
1559,38
1560,39
1561,39
1562,39
1563,39
1564,39
1565,39
1566,39
1567,39
1568,39
1569,39
1570,39
1571,39
1572,39
1573,39
1574,39
1575,39
1576,39
1577,39
1578,39
1579,39
1580,39
1581,39
1582,39
1583,39
1584,39
1585,39
1586,39
1587,39
1588,39
1589,39
1590,39
1591,39
1592,39
1593,39
1594,39
1595,39
1596,39
1597,39
1598,39
1599,39
1600,40
1601,40
1602,40
1603,40
1604,40
1605,40
1606,40
1607,40
1608,40
1609,40
1610,40
1611,40
1612,40
1613,40
1614,40
1615,40
1616,40
1617,40
1618,40
1619,40
1620,40
1621,40
1622,40
1623,40
1624,40
1625,40
1626,40
1627,40
1628,40
1629,40
1630,40
1631,40
1632,40
1633,40
1634,40
1635,40
1636,40
1637,40
1638,40
1639,40
1640,41
1641,41
1642,41
1643,41
1644,41
1645,41
1646,41
1647,41
1648,41
1649,41
1650,41
1651,41
1652,41
1653,41
1654,41
1655,41
1656,41
1657,41
1658,41
1659,41
1660,41
1661,41
1662,41
1663,41
1664,41
1665,41
1666,41
1667,41
1668,41
1669,41
1670,41
1671,41
1672,41
1673,41
1674,41
1675,41
1676,41
1677,41
1678,41
1679,41
1680,42
1681,42
1682,42
1683,42
1684,42
1685,42
1686,42
1687,42
1688,42
1689,42
1690,42
1691,42
1692,42
1693,42
1694,42
1695,42
1696,42
1697,42
1698,42
1699,42
1700,42
1701,42
1702,42
1703,42
1704,42
1705,42
1706,42
1707,42
1708,42
1709,42
1710,42
1711,42
1712,42
1713,42
1714,42
1715,42
1716,42
1717,42
1718,42
1719,42
1720,43
1721,43
1722,43
1723,43
1724,43
1725,43
1726,43
1727,43
1728,43
1729,43
1730,43
1731,43
1732,43
1733,43
1734,43
1735,43
1736,43
1737,43
1738,43
1739,43
1740,43
1741,43
1742,43
1743,43
1744,43
1745,43
1746,43
1747,43
1748,43
1749,43
1750,43
1751,43
1752,43
1753,43
1754,43
1755,43
1756,43
1757,43
1758,43
1759,43
1760,44
1761,44
1762,44
1763,44
1764,44
1765,44
1766,44
1767,44
1768,44
1769,44
1770,44
1771,44
1772,44
1773,44
1774,44
1775,44
1776,44
1777,44
1778,44
1779,44
1780,44
1781,44
1782,44
1783,44
1784,44
1785,44
1786,44
1787,44
1788,44
1789,44
1790,44
1791,44
1792,44
1793,44
1794,44
1795,44
1796,44
1797,44
1798,44
1799,44
1800,45
1801,45
1802,45
1803,45
1804,45
1805,45
1806,45
1807,45
1808,45
1809,45
1810,45
1811,45
1812,45
1813,45
1814,45
1815,45
1816,45
1817,45
1818,45
1819,45
1820,45
1821,45
1822,45
1823,45
1824,45
1825,45
1826,45
1827,45
1828,45
1829,45
1830,45
1831,45
1832,45
1833,45
1834,45
1835,45
1836,45
1837,45
1838,45
1839,45
1840,46
1841,46
1842,46
1843,46
1844,46
1845,46
1846,46
1847,46
1848,46
1849,46
1850,46
1851,46
1852,46
1853,46
1854,46
1855,46
1856,46
1857,46
1858,46
1859,46
1860,46
1861,46
1862,46
1863,46
1864,46
1865,46
1866,46
1867,46
1868,46
1869,46
1870,46
1871,46
1872,46
1873,46
1874,46
1875,46
1876,46
1877,46
1878,46
1879,46
1880,47
1881,47
1882,47
1883,47
1884,47
1885,47
1886,47
1887,47
1888,47
1889,47
1890,47
1891,47
1892,47
1893,47
1894,47
1895,47
1896,47
1897,47
1898,47
1899,47
1900,47
1901,47
1902,47
1903,47
1904,47
1905,47
1906,47
1907,47
1908,47
1909,47
1910,47
1911,47
1912,47
1913,47
1914,47
1915,47
1916,47
1917,47
1918,47
1919,47
1920,48
1921,48
1922,48
1923,48
1924,48
1925,48
1926,48
1927,48
1928,48
1929,48
1930,48
1931,48
1932,48
1933,48
1934,48
1935,48
1936,48
1937,48
1938,48
1939,48
1940,48
1941,48
1942,48
1943,48
1944,48
1945,48
1946,48
1947,48
1948,48
1949,48
1950,48
1951,48
1952,48
1953,48
1954,48
1955,48
1956,48
1957,48
1958,48
1959,48
1960,49
1961,49
1962,49
1963,49
1964,49
1965,49
1966,49
1967,49
1968,49
1969,49
1970,49
1971,49
1972,49
1973,49
1974,49
1975,49
1976,49
1977,49
1978,49
1979,49
1980,49
1981,49
1982,49
1983,49
1984,49
1985,49
1986,49
1987,49
1988,49
1989,49
1990,49
1991,49
1992,49
1993,49
1994,49
1995,49
1996,49
1997,49
1998,49
1999,49
2000,50
2001,50
2002,50
2003,50
2004,50
2005,50
2006,50
2007,50
2008,50
2009,50
2010,50
2011,50
2012,50
2013,50
2014,50
2015,50
2016,50
2017,50
2018,50
2019,50
2020,50
2021,50
2022,50
2023,50
2024,50
2025,50
2026,50
2027,50
2028,50
2029,50
2030,50
2031,50
2032,50
2033,50
2034,50
2035,50
2036,50
2037,50
2038,50
2039,50
2040,51
2041,51
2042,51
2043,51
2044,51
2045,51
2046,51
2047,51
2048,51
2049,51
2050,51
2051,51
2052,51
2053,51
2054,51
2055,51
2056,51
2057,51
2058,51
2059,51
2060,51
2061,51
2062,51
2063,51
2064,51
2065,51
2066,51
2067,51
2068,51
2069,51
2070,51
2071,51
2072,51
2073,51
2074,51
2075,51
2076,51
2077,51
2078,51
2079,51
2080,52
2081,52
2082,52
2083,52
2084,52
2085,52
2086,52
2087,52
2088,52
2089,52
2090,52
2091,52
2092,52
2093,52
2094,52
2095,52
2096,52
2097,52
2098,52
2099,52
2100,52
2101,52
2102,52
2103,52
2104,52
2105,52
2106,52
2107,52
2108,52
2109,52
2110,52
2111,52
2112,52
2113,52
2114,52
2115,52
2116,52
2117,52
2118,52
2119,52
2120,53
2121,53
2122,53
2123,53
2124,53
2125,53
2126,53
2127,53
2128,53
2129,53
2130,53
2131,53
2132,53
2133,53
2134,53
2135,53
2136,53
2137,53
2138,53
2139,53
2140,53
2141,53
2142,53
2143,53
2144,53
2145,53
2146,53
2147,53
2148,53
2149,53
2150,53
2151,53
2152,53
2153,53
2154,53
2155,53
2156,53
2157,53
2158,53
2159,53
2160,54
2161,54
2162,54
2163,54
2164,54
2165,54
2166,54
2167,54
2168,54
2169,54
2170,54
2171,54
2172,54
2173,54
2174,54
2175,54
2176,54
2177,54
2178,54
2179,54
2180,54
2181,54
2182,54
2183,54
2184,54
2185,54
2186,54
2187,54
2188,54
2189,54
2190,54
2191,54
2192,54
2193,54
2194,54
2195,54
2196,54
2197,54
2198,54
2199,54
2200,55
2201,55
2202,55
2203,55
2204,55
2205,55
2206,55
2207,55
2208,55
2209,55
2210,55
2211,55
2212,55
2213,55
2214,55
2215,55
2216,55
2217,55
2218,55
2219,55
2220,55
2221,55
2222,55
2223,55
2224,55
2225,55
2226,55
2227,55
2228,55
2229,55
2230,55
2231,55
2232,55
2233,55
2234,55
2235,55
2236,55
2237,55
2238,55
2239,55
2240,56
2241,56
2242,56
2243,56
2244,56
2245,56
2246,56
2247,56
2248,56
2249,56
2250,56
2251,56
2252,56
2253,56
2254,56
2255,56
2256,56
2257,56
2258,56
2259,56
2260,56
2261,56
2262,56
2263,56
2264,56
2265,56
2266,56
2267,56
2268,56
2269,56
2270,56
2271,56
2272,56
2273,56
2274,56
2275,56
2276,56
2277,56
2278,56
2279,56
2280,57
2281,57
2282,57
2283,57
2284,57
2285,57
2286,57
2287,57
2288,57
2289,57
2290,57
2291,57
2292,57
2293,57
2294,57
2295,57
2296,57
2297,57
2298,57
2299,57
2300,57
2301,57
2302,57
2303,57
2304,57
2305,57
2306,57
2307,57
2308,57
2309,57
2310,57
2311,57
2312,57
2313,57
2314,57
2315,57
2316,57
2317,57
2318,57
2319,57
2320,58
2321,58
2322,58
2323,58
2324,58
2325,58
2326,58
2327,58
2328,58
2329,58
2330,58
2331,58
2332,58
2333,58
2334,58
2335,58
2336,58
2337,58
2338,58
2339,58
2340,58
2341,58
2342,58
2343,58
2344,58
2345,58
2346,58
2347,58
2348,58
2349,58
2350,58
2351,58
2352,58
2353,58
2354,58
2355,58
2356,58
2357,58
2358,58
2359,58
2360,59
2361,59
2362,59
2363,59
2364,59
2365,59
2366,59
2367,59
2368,59
2369,59
2370,59
2371,59
2372,59
2373,59
2374,59
2375,59
2376,59
2377,59
2378,59
2379,59
2380,59
2381,59
2382,59
2383,59
2384,59
2385,59
2386,59
2387,59
2388,59
2389,59
2390,59
2391,59
2392,59
2393,59
2394,59
2395,59
2396,59
2397,59
2398,59
2399,59
2400,60
2401,60
2402,60
2403,60
2404,60
2405,60
2406,60
2407,60
2408,60
2409,60
2410,60
2411,60
2412,60
2413,60
2414,60
2415,60
2416,60
2417,60
2418,60
2419,60
2420,60
2421,60
2422,60
2423,60
2424,60
2425,60
2426,60
2427,60
2428,60
2429,60
2430,60
2431,60
2432,60
2433,60
2434,60
2435,60
2436,60
2437,60
2438,60
2439,60
2440,61
2441,61
2442,61
2443,61
2444,61
2445,61
2446,61
2447,61
2448,61
2449,61
2450,61
2451,61
2452,61
2453,61
2454,61
2455,61
2456,61
2457,61
2458,61
2459,61
2460,61
2461,61
2462,61
2463,61
2464,61
2465,61
2466,61
2467,61
2468,61
2469,61
2470,61
2471,61
2472,61
2473,61
2474,61
2475,61
2476,61
2477,61
2478,61
2479,61
2480,62
2481,62
2482,62
2483,62
2484,62
2485,62
2486,62
2487,62
2488,62
2489,62
2490,62
2491,62
2492,62
2493,62
2494,62
2495,62
2496,62
2497,62
2498,62
2499,62
2500,62
2501,62
2502,62
2503,62
2504,62
2505,62
2506,62
2507,62
2508,62
2509,62
2510,62
2511,62
2512,62
2513,62
2514,62
2515,62
2516,62
2517,62
2518,62
2519,62
2520,63
2521,63
2522,63
2523,63
2524,63
2525,63
2526,63
2527,63
2528,63
2529,63
2530,63
2531,63
2532,63
2533,63
2534,63
2535,63
2536,63
2537,63
2538,63
2539,63
2540,63
2541,63
2542,63
2543,63
2544,63
2545,63
2546,63
2547,63
2548,63
2549,63
2550,63
2551,63
2552,63
2553,63
2554,63
2555,63
2556,63
2557,63
2558,63
2559,63
2560,64
2561,64
2562,64
2563,64
2564,64
2565,64
2566,64
2567,64
2568,64
2569,64
2570,64
2571,64
2572,64
2573,64
2574,64
2575,64
2576,64
2577,64
2578,64
2579,64
2580,64
2581,64
2582,64
2583,64
2584,64
2585,64
2586,64
2587,64
2588,64
2589,64
2590,64
2591,64
2592,64
2593,64
2594,64
2595,64
2596,64
2597,64
2598,64
2599,64
2600,65
2601,65
2602,65
2603,65
2604,65
2605,65
2606,65
2607,65
2608,65
2609,65
2610,65
2611,65
2612,65
2613,65
2614,65
2615,65
2616,65
2617,65
2618,65
2619,65
2620,65
2621,65
2622,65
2623,65
2624,65
2625,65
2626,65
2627,65
2628,65
2629,65
2630,65
2631,65
2632,65
2633,65
2634,65
2635,65
2636,65
2637,65
2638,65
2639,65
2640,66
2641,66
2642,66
2643,66
2644,66
2645,66
2646,66
2647,66
2648,66
2649,66
2650,66
2651,66
2652,66
2653,66
2654,66
2655,66
2656,66
2657,66
2658,66
2659,66
2660,66
2661,66
2662,66
2663,66
2664,66
2665,66
2666,66
2667,66
2668,66
2669,66
2670,66
2671,66
2672,66
2673,66
2674,66
2675,66
2676,66
2677,66
2678,66
2679,66
2680,67
2681,67
2682,67
2683,67
2684,67
2685,67
2686,67
2687,67
2688,67
2689,67
2690,67
2691,67
2692,67
2693,67
2694,67
2695,67
2696,67
2697,67
2698,67
2699,67
2700,67
2701,67
2702,67
2703,67
2704,67
2705,67
2706,67
2707,67
2708,67
2709,67
2710,67
2711,67
2712,67
2713,67
2714,67
2715,67
2716,67
2717,67
2718,67
2719,67
2720,68
2721,68
2722,68
2723,68
2724,68
2725,68
2726,68
2727,68
2728,68
2729,68
2730,68
2731,68
2732,68
2733,68
2734,68
2735,68
2736,68
2737,68
2738,68
2739,68
2740,68
2741,68
2742,68
2743,68
2744,68
2745,68
2746,68
2747,68
2748,68
2749,68
2750,68
2751,68
2752,68
2753,68
2754,68
2755,68
2756,68
2757,68
2758,68
2759,68
2760,69
2761,69
2762,69
2763,69
2764,69
2765,69
2766,69
2767,69
2768,69
2769,69
2770,69
2771,69
2772,69
2773,69
2774,69
2775,69
2776,69
2777,69
2778,69
2779,69
2780,69
2781,69
2782,69
2783,69
2784,69
2785,69
2786,69
2787,69
2788,69
2789,69
2790,69
2791,69
2792,69
2793,69
2794,69
2795,69
2796,69
2797,69
2798,69
2799,69
2800,70
2801,70
2802,70
2803,70
2804,70
2805,70
2806,70
2807,70
2808,70
2809,70
2810,70
2811,70
2812,70
2813,70
2814,70
2815,70
2816,70
2817,70
2818,70
2819,70
2820,70
2821,70
2822,70
2823,70
2824,70
2825,70
2826,70
2827,70
2828,70
2829,70
2830,70
2831,70
2832,70
2833,70
2834,70
2835,70
2836,70
2837,70
2838,70
2839,70
2840,71
2841,71
2842,71
2843,71
2844,71
2845,71
2846,71
2847,71
2848,71
2849,71
2850,71
2851,71
2852,71
2853,71
2854,71
2855,71
2856,71
2857,71
2858,71
2859,71
2860,71
2861,71
2862,71
2863,71
2864,71
2865,71
2866,71
2867,71
2868,71
2869,71
2870,71
2871,71
2872,71
2873,71
2874,71
2875,71
2876,71
2877,71
2878,71
2879,71
2880,72
2881,72
2882,72
2883,72
2884,72
2885,72
2886,72
2887,72
2888,72
2889,72
2890,72
2891,72
2892,72
2893,72
2894,72
2895,72
2896,72
2897,72
2898,72
2899,72
2900,72
2901,72
2902,72
2903,72
2904,72
2905,72
2906,72
2907,72
2908,72
2909,72
2910,72
2911,72
2912,72
2913,72
2914,72
2915,72
2916,72
2917,72
2918,72
2919,72
2920,73
2921,73
2922,73
2923,73
2924,73
2925,73
2926,73
2927,73
2928,73
2929,73
2930,73
2931,73
2932,73
2933,73
2934,73
2935,73
2936,73
2937,73
2938,73
2939,73
2940,73
2941,73
2942,73
2943,73
2944,73
2945,73
2946,73
2947,73
2948,73
2949,73
2950,73
2951,73
2952,73
2953,73
2954,73
2955,73
2956,73
2957,73
2958,73
2959,73
2960,74
2961,74
2962,74
2963,74
2964,74
2965,74
2966,74
2967,74
2968,74
2969,74
2970,74
2971,74
2972,74
2973,74
2974,74
2975,74
2976,74
2977,74
2978,74
2979,74
2980,74
2981,74
2982,74
2983,74
2984,74
2985,74
2986,74
2987,74
2988,74
2989,74
2990,74
2991,74
2992,74
2993,74
2994,74
2995,74
2996,74
2997,74
2998,74
2999,74
3000,75
3001,75
3002,75
3003,75
3004,75
3005,75
3006,75
3007,75
3008,75
3009,75
3010,75
3011,75
3012,75
3013,75
3014,75
3015,75
3016,75
3017,75
3018,75
3019,75
3020,75
3021,75
3022,75
3023,75
3024,75
3025,75
3026,75
3027,75
3028,75
3029,75
3030,75
3031,75
3032,75
3033,75
3034,75
3035,75
3036,75
3037,75
3038,75
3039,75
3040,76
3041,76
3042,76
3043,76
3044,76
3045,76
3046,76
3047,76
3048,76
3049,76
3050,76
3051,76
3052,76
3053,76
3054,76
3055,76
3056,76
3057,76
3058,76
3059,76
3060,76
3061,76
3062,76
3063,76
3064,76
3065,76
3066,76
3067,76
3068,76
3069,76
3070,76
3071,76
3072,76
3073,76
3074,76
3075,76
3076,76
3077,76
3078,76
3079,76
3080,77
3081,77
3082,77
3083,77
3084,77
3085,77
3086,77
3087,77
3088,77
3089,77
3090,77
3091,77
3092,77
3093,77
3094,77
3095,77
3096,77
3097,77
3098,77
3099,77
3100,77
3101,77
3102,77
3103,77
3104,77
3105,77
3106,77
3107,77
3108,77
3109,77
3110,77
3111,77
3112,77
3113,77
3114,77
3115,77
3116,77
3117,77
3118,77
3119,77
