0,0
1,0
2,0
3,0
4,0
5,0
6,0
7,0
8,0
9,0
10,0
11,0
12,0
13,0
14,0
15,0
16,0
17,0
18,0
19,0
20,0
21,0
22,0
23,0
24,0
25,0
26,0
27,0
28,0
29,0
30,0
31,0
32,0
33,0
34,0
35,0
36,0
37,0
38,1
39,1
40,1
41,1
42,1
43,1
44,1
45,1
46,1
47,1
48,1
49,1
50,1
51,1
52,1
53,1
54,1
55,1
56,1
57,1
58,1
59,1
60,1
61,1
62,1
63,1
64,1
65,1
66,1
67,1
68,1
69,1
70,1
71,1
72,1
73,1
74,1
75,1
76,2
77,2
78,2
79,2
80,2
81,2
82,2
83,2
84,2
85,2
86,2
87,2
88,2
89,2
90,2
91,2
92,2
93,2
94,2
95,2
96,2
97,2
98,2
99,2
100,2
101,2
102,2
103,2
104,2
105,2
106,2
107,2
108,2
109,2
110,2
111,2
112,2
113,2
114,3
115,3
116,3
117,3
118,3
119,3
120,3
121,3
122,3
123,3
124,3
125,3
126,3
127,3
128,3
129,3
130,3
131,3
132,3
133,3
134,3
135,3
136,3
137,3
138,3
139,3
140,3
141,3
142,3
143,3
144,3
145,3
146,3
147,3
148,3
149,3
150,3
151,3
152,4
153,4
154,4
155,4
156,4
157,4
158,4
159,4
160,4
161,4
162,4
163,4
164,4
165,4
166,4
167,4
168,4
169,4
170,4
171,4
172,4
173,4
174,4
175,4
176,4
177,4
178,4
179,4
180,4
181,4
182,4
183,4
184,4
185,4
186,4
187,4
188,4
189,4
190,5
191,5
192,5
193,5
194,5
195,5
196,5
197,5
198,5
199,5
200,5
201,5
202,5
203,5
204,5
205,5
206,5
207,5
208,5
209,5
210,5
211,5
212,5
213,5
214,5
215,5
216,5
217,5
218,5
219,5
220,5
221,5
222,5
223,5
224,5
225,5
226,5
227,5
228,6
229,6
230,6
231,6
232,6
233,6
234,6
235,6
236,6
237,6
238,6
239,6
240,6
241,6
242,6
243,6
244,6
245,6
246,6
247,6
248,6
249,6
250,6
251,6
252,6
253,6
254,6
255,6
256,6
257,6
258,6
259,6
260,6
261,6
262,6
263,6
264,6
265,6
266,7
267,7
268,7
269,7
270,7
271,7
272,7
273,7
274,7
275,7
276,7
277,7
278,7
279,7
280,7
281,7
282,7
283,7
284,7
285,7
286,7
287,7
288,7
289,7
290,7
291,7
292,7
293,7
294,7
295,7
296,7
297,7
298,7
299,7
300,7
301,7
302,7
303,7
304,8
305,8
306,8
307,8
308,8
309,8
310,8
311,8
312,8
313,8
314,8
315,8
316,8
317,8
318,8
319,8
320,8
321,8
322,8
323,8
324,8
325,8
326,8
327,8
328,8
329,8
330,8
331,8
332,8
333,8
334,8
335,8
336,8
337,8
338,8
339,8
340,8
341,8
342,9
343,9
344,9
345,9
346,9
347,9
348,9
349,9
350,9
351,9
352,9
353,9
354,9
355,9
356,9
357,9
358,9
359,9
360,9
361,9
362,9
363,9
364,9
365,9
366,9
367,9
368,9
369,9
370,9
371,9
372,9
373,9
374,9
375,9
376,9
377,9
378,9
379,9
380,10
381,10
382,10
383,10
384,10
385,10
386,10
387,10
388,10
389,10
390,10
391,10
392,10
393,10
394,10
395,10
396,10
397,10
398,10
399,10
400,10
401,10
402,10
403,10
404,10
405,10
406,10
407,10
408,10
409,10
410,10
411,10
412,10
413,10
414,10
415,10
416,10
417,10
418,11
419,11
420,11
421,11
422,11
423,11
424,11
425,11
426,11
427,11
428,11
429,11
430,11
431,11
432,11
433,11
434,11
435,11
436,11
437,11
438,11
439,11
440,11
441,11
442,11
443,11
444,11
445,11
446,11
447,11
448,11
449,11
450,11
451,11
452,11
453,11
454,11
455,11
456,12
457,12
458,12
459,12
460,12
461,12
462,12
463,12
464,12
465,12
466,12
467,12
468,12
469,12
470,12
471,12
472,12
473,12
474,12
475,12
476,12
477,12
478,12
479,12
480,12
481,12
482,12
483,12
484,12
485,12
486,12
487,12
488,12
489,12
490,12
491,12
492,12
493,12
494,13
495,13
496,13
497,13
498,13
499,13
500,13
501,13
502,13
503,13
504,13
505,13
506,13
507,13
508,13
509,13
510,13
511,13
512,13
513,13
514,13
515,13
516,13
517,13
518,13
519,13
520,13
521,13
522,13
523,13
524,13
525,13
526,13
527,13
528,13
529,13
530,13
531,13
532,14
533,14
534,14
535,14
536,14
537,14
538,14
539,14
540,14
541,14
542,14
543,14
544,14
545,14
546,14
547,14
548,14
549,14
550,14
551,14
552,14
553,14
554,14
555,14
556,14
557,14
558,14
559,14
560,14
561,14
562,14
563,14
564,14
565,14
566,14
567,14
568,15
569,15
570,15
571,15
572,15
573,15
574,15
575,15
576,15
577,15
578,15
579,15
580,15
581,15
582,15
583,15
584,15
585,15
586,15
587,15
588,15
589,15
590,15
591,15
592,15
593,15
594,15
595,15
596,15
597,15
598,15
599,15
600,15
601,15
602,15
603,15
604,16
605,16
606,16
607,16
608,16
609,16
610,16
611,16
612,16
613,16
614,16
615,16
616,16
617,16
618,16
619,16
620,16
621,16
622,16
623,16
624,16
625,16
626,16
627,16
628,16
629,16
630,16
631,16
632,16
633,16
634,16
635,16
636,16
637,16
638,16
639,16
640,17
641,17
642,17
643,17
644,17
645,17
646,17
647,17
648,17
649,17
650,17
651,17
652,17
653,17
654,17
655,17
656,17
657,17
658,17
659,17
660,17
661,17
662,17
663,17
664,17
665,17
666,17
667,17
668,17
669,17
670,17
671,17
672,17
673,17
674,17
675,17
676,18
677,18
678,18
679,18
680,18
681,18
682,18
683,18
684,18
685,18
686,18
687,18
688,18
689,18
690,18
691,18
692,18
693,18
694,18
695,18
696,18
697,18
698,18
699,18
700,18
701,18
702,18
703,18
704,18
705,18
706,18
707,18
708,18
709,18
710,18
711,18
712,19
713,19
714,19
715,19
716,19
717,19
718,19
719,19
720,19
721,19
722,19
723,19
724,19
725,19
726,19
727,19
728,19
729,19
730,19
731,19
732,19
733,19
734,19
735,19
736,19
737,19
738,19
739,19
740,19
741,19
742,19
743,19
744,19
745,19
746,19
747,19
748,20
749,20
750,20
751,20
752,20
753,20
754,20
755,20
756,20
757,20
758,20
759,20
760,20
761,20
762,20
763,20
764,20
765,20
766,20
767,20
768,20
769,20
770,20
771,20
772,20
773,20
774,20
775,20
776,20
777,20
778,20
779,20
780,20
781,20
782,20
783,20
784,20
785,20
786,21
787,21
788,21
789,21
790,21
791,21
792,21
793,21
794,21
795,21
796,21
797,21
798,21
799,21
800,21
801,21
802,21
803,21
804,21
805,21
806,21
807,21
808,21
809,21
810,21
811,21
812,21
813,21
814,21
815,21
816,21
817,21
818,21
819,21
820,21
821,21
822,21
823,21
824,22
825,22
826,22
827,22
828,22
829,22
830,22
831,22
832,22
833,22
834,22
835,22
836,22
837,22
838,22
839,22
840,22
841,22
842,22
843,22
844,22
845,22
846,22
847,22
848,22
849,22
850,22
851,22
852,22
853,22
854,22
855,22
856,22
857,22
858,22
859,22
860,22
861,22
862,23
863,23
864,23
865,23
866,23
867,23
868,23
869,23
870,23
871,23
872,23
873,23
874,23
875,23
876,23
877,23
878,23
879,23
880,23
881,23
882,23
883,23
884,23
885,23
886,23
887,23
888,23
889,23
890,23
891,23
892,23
893,23
894,23
895,23
896,23
897,23
898,23
899,23
900,24
901,24
902,24
903,24
904,24
905,24
906,24
907,24
908,24
909,24
910,24
911,24
912,24
913,24
914,24
915,24
916,24
917,24
918,24
919,24
920,24
921,24
922,24
923,24
924,24
925,24
926,24
927,24
928,24
929,24
930,24
931,24
932,24
933,24
934,24
935,24
936,24
937,24
938,25
939,25
940,25
941,25
942,25
943,25
944,25
945,25
946,25
947,25
948,25
949,25
950,25
951,25
952,25
953,25
954,25
955,25
956,25
957,25
958,25
959,25
960,25
961,25
962,25
963,25
964,25
965,25
966,25
967,25
968,25
969,25
970,25
971,25
972,25
973,25
974,25
975,25
976,26
977,26
978,26
979,26
980,26
981,26
982,26
983,26
984,26
985,26
986,26
987,26
988,26
989,26
990,26
991,26
992,26
993,26
994,26
995,26
996,26
997,26
998,26
999,26
1000,26
1001,26
1002,26
1003,26
1004,26
1005,26
1006,26
1007,26
1008,26
1009,26
1010,26
1011,26
1012,26
1013,26
1014,27
1015,27
1016,27
1017,27
1018,27
1019,27
1020,27
1021,27
1022,27
1023,27
1024,27
1025,27
1026,27
1027,27
1028,27
1029,27
1030,27
1031,27
1032,27
1033,27
1034,27
1035,27
1036,27
1037,27
1038,27
1039,27
1040,27
1041,27
1042,27
1043,27
1044,27
1045,27
1046,27
1047,27
1048,27
1049,27
1050,27
1051,27
1052,28
1053,28
1054,28
1055,28
1056,28
1057,28
1058,28
1059,28
1060,28
1061,28
1062,28
1063,28
1064,28
1065,28
1066,28
1067,28
1068,28
1069,28
1070,28
1071,28
1072,28
1073,28
1074,28
1075,28
1076,28
1077,28
1078,28
1079,28
1080,28
1081,28
1082,28
1083,28
1084,28
1085,28
1086,28
1087,28
1088,28
1089,28
1090,29
1091,29
1092,29
1093,29
1094,29
1095,29
1096,29
1097,29
1098,29
1099,29
1100,29
1101,29
1102,29
1103,29
1104,29
1105,29
1106,29
1107,29
1108,29
1109,29
1110,29
1111,29
1112,29
1113,29
1114,29
1115,29
1116,29
1117,29
1118,29
1119,29
1120,29
1121,29
1122,29
1123,29
1124,29
1125,29
1126,29
1127,29
1128,30
1129,30
1130,30
1131,30
1132,30
1133,30
1134,30
1135,30
1136,30
1137,30
1138,30
1139,30
1140,30
1141,30
1142,30
1143,30
1144,30
1145,30
1146,30
1147,30
1148,30
1149,30
1150,30
1151,30
1152,30
1153,30
1154,30
1155,30
1156,30
1157,30
1158,30
1159,30
1160,30
1161,30
1162,30
1163,30
1164,30
1165,30
1166,31
1167,31
1168,31
1169,31
1170,31
1171,31
1172,31
1173,31
1174,31
1175,31
1176,31
1177,31
1178,31
1179,31
1180,31
1181,31
1182,31
1183,31
1184,31
1185,31
1186,31
1187,31
1188,31
1189,31
1190,31
1191,31
1192,31
1193,31
1194,31
1195,31
1196,31
1197,31
1198,31
1199,31
1200,31
1201,31
1202,31
1203,31
1204,32
1205,32
1206,32
1207,32
1208,32
1209,32
1210,32
1211,32
1212,32
1213,32
1214,32
1215,32
1216,32
1217,32
1218,32
1219,32
1220,32
1221,32
1222,32
1223,32
1224,32
1225,32
1226,32
1227,32
1228,32
1229,32
1230,32
1231,32
1232,32
1233,32
1234,32
1235,32
1236,32
1237,32
1238,32
1239,32
1240,32
1241,32
1242,33
1243,33
1244,33
1245,33
1246,33
1247,33
1248,33
1249,33
1250,33
1251,33
1252,33
1253,33
1254,33
1255,33
1256,33
1257,33
1258,33
1259,33
1260,33
1261,33
1262,33
1263,33
1264,33
1265,33
1266,33
1267,33
1268,33
1269,33
1270,33
1271,33
1272,33
1273,33
1274,33
1275,33
1276,33
1277,33
1278,33
1279,33
1280,34
1281,34
1282,34
1283,34
1284,34
1285,34
1286,34
1287,34
1288,34
1289,34
1290,34
1291,34
1292,34
1293,34
1294,34
1295,34
1296,34
1297,34
1298,34
1299,34
1300,34
1301,34
1302,34
1303,34
1304,34
1305,34
1306,34
1307,34
1308,34
1309,34
1310,34
1311,34
1312,34
1313,34
1314,34
1315,34
1316,35
1317,35
1318,35
1319,35
1320,35
1321,35
1322,35
1323,35
1324,35
1325,35
1326,35
1327,35
1328,35
1329,35
1330,35
1331,35
1332,35
1333,35
1334,35
1335,35
1336,35
1337,35
1338,35
1339,35
1340,35
1341,35
1342,35
1343,35
1344,35
1345,35
1346,35
1347,35
1348,35
1349,35
1350,35
1351,35
1352,36
1353,36
1354,36
1355,36
1356,36
1357,36
1358,36
1359,36
1360,36
1361,36
1362,36
1363,36
1364,36
1365,36
1366,36
1367,36
1368,36
1369,36
1370,36
1371,36
1372,36
1373,36
1374,36
1375,36
1376,36
1377,36
1378,36
1379,36
1380,36
1381,36
1382,36
1383,36
1384,36
1385,36
1386,36
1387,36
1388,37
1389,37
1390,37
1391,37
1392,37
1393,37
1394,37
1395,37
1396,37
1397,37
1398,37
1399,37
1400,37
1401,37
1402,37
1403,37
1404,37
1405,37
1406,37
1407,37
1408,37
1409,37
1410,37
1411,37
1412,37
1413,37
1414,37
1415,37
1416,37
1417,37
1418,37
1419,37
1420,37
1421,37
1422,37
1423,37
1424,38
1425,38
1426,38
1427,38
1428,38
1429,38
1430,38
1431,38
1432,38
1433,38
1434,38
1435,38
1436,38
1437,38
1438,38
1439,38
1440,38
1441,38
1442,38
1443,38
1444,38
1445,38
1446,38
1447,38
1448,38
1449,38
1450,38
1451,38
1452,38
1453,38
1454,38
1455,38
1456,38
1457,38
1458,38
1459,38
1460,39
1461,39
1462,39
1463,39
1464,39
1465,39
1466,39
1467,39
1468,39
1469,39
1470,39
1471,39
1472,39
1473,39
1474,39
1475,39
1476,39
1477,39
1478,39
1479,39
1480,39
1481,39
1482,39
1483,39
1484,39
1485,39
1486,39
1487,39
1488,39
1489,39
1490,39
1491,39
1492,39
1493,39
1494,39
1495,39
1496,40
1497,40
1498,40
1499,40
1500,40
1501,40
1502,40
1503,40
1504,40
1505,40
1506,40
1507,40
1508,40
1509,40
1510,40
1511,40
1512,40
1513,40
1514,40
1515,40
1516,40
1517,40
1518,40
1519,40
1520,40
1521,40
1522,40
1523,40
1524,40
1525,40
1526,40
1527,40
1528,40
1529,40
1530,40
1531,40
1532,40
1533,40
1534,41
1535,41
1536,41
1537,41
1538,41
1539,41
1540,41
1541,41
1542,41
1543,41
1544,41
1545,41
1546,41
1547,41
1548,41
1549,41
1550,41
1551,41
1552,41
1553,41
1554,41
1555,41
1556,41
1557,41
1558,41
1559,41
1560,41
1561,41
1562,41
1563,41
1564,41
1565,41
1566,41
1567,41
1568,41
1569,41
1570,41
1571,41
1572,42
1573,42
1574,42
1575,42
1576,42
1577,42
1578,42
1579,42
1580,42
1581,42
1582,42
1583,42
1584,42
1585,42
1586,42
1587,42
1588,42
1589,42
1590,42
1591,42
1592,42
1593,42
1594,42
1595,42
1596,42
1597,42
1598,42
1599,42
1600,42
1601,42
1602,42
1603,42
1604,42
1605,42
1606,42
1607,42
1608,42
1609,42
1610,43
1611,43
1612,43
1613,43
1614,43
1615,43
1616,43
1617,43
1618,43
1619,43
1620,43
1621,43
1622,43
1623,43
1624,43
1625,43
1626,43
1627,43
1628,43
1629,43
1630,43
1631,43
1632,43
1633,43
1634,43
1635,43
1636,43
1637,43
1638,43
1639,43
1640,43
1641,43
1642,43
1643,43
1644,43
1645,43
1646,43
1647,43
1648,44
1649,44
1650,44
1651,44
1652,44
1653,44
1654,44
1655,44
1656,44
1657,44
1658,44
1659,44
1660,44
1661,44
1662,44
1663,44
1664,44
1665,44
1666,44
1667,44
1668,44
1669,44
1670,44
1671,44
1672,44
1673,44
1674,44
1675,44
1676,44
1677,44
1678,44
1679,44
1680,44
1681,44
1682,44
1683,44
1684,44
1685,44
1686,45
1687,45
1688,45
1689,45
1690,45
1691,45
1692,45
1693,45
1694,45
1695,45
1696,45
1697,45
1698,45
1699,45
1700,45
1701,45
1702,45
1703,45
1704,45
1705,45
1706,45
1707,45
1708,45
1709,45
1710,45
1711,45
1712,45
1713,45
1714,45
1715,45
1716,45
1717,45
1718,45
1719,45
1720,45
1721,45
1722,45
1723,45
1724,46
1725,46
1726,46
1727,46
1728,46
1729,46
1730,46
1731,46
1732,46
1733,46
1734,46
1735,46
1736,46
1737,46
1738,46
1739,46
1740,46
1741,46
1742,46
1743,46
1744,46
1745,46
1746,46
1747,46
1748,46
1749,46
1750,46
1751,46
1752,46
1753,46
1754,46
1755,46
1756,46
1757,46
1758,46
1759,46
1760,46
1761,46
1762,47
1763,47
1764,47
1765,47
1766,47
1767,47
1768,47
1769,47
1770,47
1771,47
1772,47
1773,47
1774,47
1775,47
1776,47
1777,47
1778,47
1779,47
1780,47
1781,47
1782,47
1783,47
1784,47
1785,47
1786,47
1787,47
1788,47
1789,47
1790,47
1791,47
1792,47
1793,47
1794,47
1795,47
1796,47
1797,47
1798,47
1799,47
1800,48
1801,48
1802,48
1803,48
1804,48
1805,48
1806,48
1807,48
1808,48
1809,48
1810,48
1811,48
1812,48
1813,48
1814,48
1815,48
1816,48
1817,48
1818,48
1819,48
1820,48
1821,48
1822,48
1823,48
1824,48
1825,48
1826,48
1827,48
1828,48
1829,48
1830,48
1831,48
1832,48
1833,48
1834,48
1835,48
1836,48
1837,48
1838,49
1839,49
1840,49
1841,49
1842,49
1843,49
1844,49
1845,49
1846,49
1847,49
1848,49
1849,49
1850,49
1851,49
1852,49
1853,49
1854,49
1855,49
1856,49
1857,49
1858,49
1859,49
1860,49
1861,49
1862,49
1863,49
1864,49
1865,49
1866,49
1867,49
1868,49
1869,49
1870,49
1871,49
1872,49
1873,49
1874,49
1875,49
1876,50
1877,50
1878,50
1879,50
1880,50
1881,50
1882,50
1883,50
1884,50
1885,50
1886,50
1887,50
1888,50
1889,50
1890,50
1891,50
1892,50
1893,50
1894,50
1895,50
1896,50
1897,50
1898,50
1899,50
1900,50
1901,50
1902,50
1903,50
1904,50
1905,50
1906,50
1907,50
1908,50
1909,50
1910,50
1911,50
1912,50
1913,50
1914,51
1915,51
1916,51
1917,51
1918,51
1919,51
1920,51
1921,51
1922,51
1923,51
1924,51
1925,51
1926,51
1927,51
1928,51
1929,51
1930,51
1931,51
1932,51
1933,51
1934,51
1935,51
1936,51
1937,51
1938,51
1939,51
1940,51
1941,51
1942,51
1943,51
1944,51
1945,51
1946,51
1947,51
1948,51
1949,51
1950,51
1951,51
1952,52
1953,52
1954,52
1955,52
1956,52
1957,52
1958,52
1959,52
1960,52
1961,52
1962,52
1963,52
1964,52
1965,52
1966,52
1967,52
1968,52
1969,52
1970,52
1971,52
1972,52
1973,52
1974,52
1975,52
1976,52
1977,52
1978,52
1979,52
1980,52
1981,52
1982,52
1983,52
1984,52
1985,52
1986,52
1987,52
1988,52
1989,52
1990,53
1991,53
1992,53
1993,53
1994,53
1995,53
1996,53
1997,53
1998,53
1999,53
2000,53
2001,53
2002,53
2003,53
2004,53
2005,53
2006,53
2007,53
2008,53
2009,53
2010,53
2011,53
2012,53
2013,53
2014,53
2015,53
2016,53
2017,53
2018,53
2019,53
2020,53
2021,53
2022,53
2023,53
2024,53
2025,53
2026,53
2027,53
2028,54
2029,54
2030,54
2031,54
2032,54
2033,54
2034,54
2035,54
2036,54
2037,54
2038,54
2039,54
2040,54
2041,54
2042,54
2043,54
2044,54
2045,54
2046,54
2047,54
2048,54
2049,54
2050,54
2051,54
2052,54
2053,54
2054,54
2055,54
2056,54
2057,54
2058,54
2059,54
2060,54
2061,54
2062,54
2063,54
2064,55
2065,55
2066,55
2067,55
2068,55
2069,55
2070,55
2071,55
2072,55
2073,55
2074,55
2075,55
2076,55
2077,55
2078,55
2079,55
2080,55
2081,55
2082,55
2083,55
2084,55
2085,55
2086,55
2087,55
2088,55
2089,55
2090,55
2091,55
2092,55
2093,55
2094,55
2095,55
2096,55
2097,55
2098,55
2099,55
2100,56
2101,56
2102,56
2103,56
2104,56
2105,56
2106,56
2107,56
2108,56
2109,56
2110,56
2111,56
2112,56
2113,56
2114,56
2115,56
2116,56
2117,56
2118,56
2119,56
2120,56
2121,56
2122,56
2123,56
2124,56
2125,56
2126,56
2127,56
2128,56
2129,56
2130,56
2131,56
2132,56
2133,56
2134,56
2135,56
2136,57
2137,57
2138,57
2139,57
2140,57
2141,57
2142,57
2143,57
2144,57
2145,57
2146,57
2147,57
2148,57
2149,57
2150,57
2151,57
2152,57
2153,57
2154,57
2155,57
2156,57
2157,57
2158,57
2159,57
2160,57
2161,57
2162,57
2163,57
2164,57
2165,57
2166,57
2167,57
2168,57
2169,57
2170,57
2171,57
2172,58
2173,58
2174,58
2175,58
2176,58
2177,58
2178,58
2179,58
2180,58
2181,58
2182,58
2183,58
2184,58
2185,58
2186,58
2187,58
2188,58
2189,58
2190,58
2191,58
2192,58
2193,58
2194,58
2195,58
2196,58
2197,58
2198,58
2199,58
2200,58
2201,58
2202,58
2203,58
2204,58
2205,58
2206,58
2207,58
2208,59
2209,59
2210,59
2211,59
2212,59
2213,59
2214,59
2215,59
2216,59
2217,59
2218,59
2219,59
2220,59
2221,59
2222,59
2223,59
2224,59
2225,59
2226,59
2227,59
2228,59
2229,59
2230,59
2231,59
2232,59
2233,59
2234,59
2235,59
2236,59
2237,59
2238,59
2239,59
2240,59
2241,59
2242,59
2243,59
2244,60
2245,60
2246,60
2247,60
2248,60
2249,60
2250,60
2251,60
2252,60
2253,60
2254,60
2255,60
2256,60
2257,60
2258,60
2259,60
2260,60
2261,60
2262,60
2263,60
2264,60
2265,60
2266,60
2267,60
2268,60
2269,60
2270,60
2271,60
2272,60
2273,60
2274,60
2275,60
2276,60
2277,60
2278,60
2279,60
2280,60
2281,60
2282,61
2283,61
2284,61
2285,61
2286,61
2287,61
2288,61
2289,61
2290,61
2291,61
2292,61
2293,61
2294,61
2295,61
2296,61
2297,61
2298,61
2299,61
2300,61
2301,61
2302,61
2303,61
2304,61
2305,61
2306,61
2307,61
2308,61
2309,61
2310,61
2311,61
2312,61
2313,61
2314,61
2315,61
2316,61
2317,61
2318,61
2319,61
2320,62
2321,62
2322,62
2323,62
2324,62
2325,62
2326,62
2327,62
2328,62
2329,62
2330,62
2331,62
2332,62
2333,62
2334,62
2335,62
2336,62
2337,62
2338,62
2339,62
2340,62
2341,62
2342,62
2343,62
2344,62
2345,62
2346,62
2347,62
2348,62
2349,62
2350,62
2351,62
2352,62
2353,62
2354,62
2355,62
2356,62
2357,62
2358,63
2359,63
2360,63
2361,63
2362,63
2363,63
2364,63
2365,63
2366,63
2367,63
2368,63
2369,63
2370,63
2371,63
2372,63
2373,63
2374,63
2375,63
2376,63
2377,63
2378,63
2379,63
2380,63
2381,63
2382,63
2383,63
2384,63
2385,63
2386,63
2387,63
2388,63
2389,63
2390,63
2391,63
2392,63
2393,63
2394,63
2395,63
2396,64
2397,64
2398,64
2399,64
2400,64
2401,64
2402,64
2403,64
2404,64
2405,64
2406,64
2407,64
2408,64
2409,64
2410,64
2411,64
2412,64
2413,64
2414,64
2415,64
2416,64
2417,64
2418,64
2419,64
2420,64
2421,64
2422,64
2423,64
2424,64
2425,64
2426,64
2427,64
2428,64
2429,64
2430,64
2431,64
2432,64
2433,64
2434,65
2435,65
2436,65
2437,65
2438,65
2439,65
2440,65
2441,65
2442,65
2443,65
2444,65
2445,65
2446,65
2447,65
2448,65
2449,65
2450,65
2451,65
2452,65
2453,65
2454,65
2455,65
2456,65
2457,65
2458,65
2459,65
2460,65
2461,65
2462,65
2463,65
2464,65
2465,65
2466,65
2467,65
2468,65
2469,65
2470,65
2471,65
2472,66
2473,66
2474,66
2475,66
2476,66
2477,66
2478,66
2479,66
2480,66
2481,66
2482,66
2483,66
2484,66
2485,66
2486,66
2487,66
2488,66
2489,66
2490,66
2491,66
2492,66
2493,66
2494,66
2495,66
2496,66
2497,66
2498,66
2499,66
2500,66
2501,66
2502,66
2503,66
2504,66
2505,66
2506,66
2507,66
2508,66
2509,66
2510,67
2511,67
2512,67
2513,67
2514,67
2515,67
2516,67
2517,67
2518,67
2519,67
2520,67
2521,67
2522,67
2523,67
2524,67
2525,67
2526,67
2527,67
2528,67
2529,67
2530,67
2531,67
2532,67
2533,67
2534,67
2535,67
2536,67
2537,67
2538,67
2539,67
2540,67
2541,67
2542,67
2543,67
2544,67
2545,67
2546,67
2547,67
2548,68
2549,68
2550,68
2551,68
2552,68
2553,68
2554,68
2555,68
2556,68
2557,68
2558,68
2559,68
2560,68
2561,68
2562,68
2563,68
2564,68
2565,68
2566,68
2567,68
2568,68
2569,68
2570,68
2571,68
2572,68
2573,68
2574,68
2575,68
2576,68
2577,68
2578,68
2579,68
2580,68
2581,68
2582,68
2583,68
2584,68
2585,68
2586,69
2587,69
2588,69
2589,69
2590,69
2591,69
2592,69
2593,69
2594,69
2595,69
2596,69
2597,69
2598,69
2599,69
2600,69
2601,69
2602,69
2603,69
2604,69
2605,69
2606,69
2607,69
2608,69
2609,69
2610,69
2611,69
2612,69
2613,69
2614,69
2615,69
2616,69
2617,69
2618,69
2619,69
2620,69
2621,69
2622,69
2623,69
2624,70
2625,70
2626,70
2627,70
2628,70
2629,70
2630,70
2631,70
2632,70
2633,70
2634,70
2635,70
2636,70
2637,70
2638,70
2639,70
2640,70
2641,70
2642,70
2643,70
2644,70
2645,70
2646,70
2647,70
2648,70
2649,70
2650,70
2651,70
2652,70
2653,70
2654,70
2655,70
2656,70
2657,70
2658,70
2659,70
2660,70
2661,70
2662,71
2663,71
2664,71
2665,71
2666,71
2667,71
2668,71
2669,71
2670,71
2671,71
2672,71
2673,71
2674,71
2675,71
2676,71
2677,71
2678,71
2679,71
2680,71
2681,71
2682,71
2683,71
2684,71
2685,71
2686,71
2687,71
2688,71
2689,71
2690,71
2691,71
2692,71
2693,71
2694,71
2695,71
2696,71
2697,71
2698,71
2699,71
2700,72
2701,72
2702,72
2703,72
2704,72
2705,72
2706,72
2707,72
2708,72
2709,72
2710,72
2711,72
2712,72
2713,72
2714,72
2715,72
2716,72
2717,72
2718,72
2719,72
2720,72
2721,72
2722,72
2723,72
2724,72
2725,72
2726,72
2727,72
2728,72
2729,72
2730,72
2731,72
2732,72
2733,72
2734,72
2735,72
2736,72
2737,72
2738,73
2739,73
2740,73
2741,73
2742,73
2743,73
2744,73
2745,73
2746,73
2747,73
2748,73
2749,73
2750,73
2751,73
2752,73
2753,73
2754,73
2755,73
2756,73
2757,73
2758,73
2759,73
2760,73
2761,73
2762,73
2763,73
2764,73
2765,73
2766,73
2767,73
2768,73
2769,73
2770,73
2771,73
2772,73
2773,73
2774,73
2775,73
2776,74
2777,74
2778,74
2779,74
2780,74
2781,74
2782,74
2783,74
2784,74
2785,74
2786,74
2787,74
2788,74
2789,74
2790,74
2791,74
2792,74
2793,74
2794,74
2795,74
2796,74
2797,74
2798,74
2799,74
2800,74
2801,74
2802,74
2803,74
2804,74
2805,74
2806,74
2807,74
2808,74
2809,74
2810,74
2811,74
2812,75
2813,75
2814,75
2815,75
2816,75
2817,75
2818,75
2819,75
2820,75
2821,75
2822,75
2823,75
2824,75
2825,75
2826,75
2827,75
2828,75
2829,75
2830,75
2831,75
2832,75
2833,75
2834,75
2835,75
2836,75
2837,75
2838,75
2839,75
2840,75
2841,75
2842,75
2843,75
2844,75
2845,75
2846,75
2847,75
2848,76
2849,76
2850,76
2851,76
2852,76
2853,76
2854,76
2855,76
2856,76
2857,76
2858,76
2859,76
2860,76
2861,76
2862,76
2863,76
2864,76
2865,76
2866,76
2867,76
2868,76
2869,76
2870,76
2871,76
2872,76
2873,76
2874,76
2875,76
2876,76
2877,76
2878,76
2879,76
2880,76
2881,76
2882,76
2883,76
2884,77
2885,77
2886,77
2887,77
2888,77
2889,77
2890,77
2891,77
2892,77
2893,77
2894,77
2895,77
2896,77
2897,77
2898,77
2899,77
2900,77
2901,77
2902,77
2903,77
2904,77
2905,77
2906,77
2907,77
2908,77
2909,77
2910,77
2911,77
2912,77
2913,77
2914,77
2915,77
2916,77
2917,77
2918,77
2919,77
2920,78
2921,78
2922,78
2923,78
2924,78
2925,78
2926,78
2927,78
2928,78
2929,78
2930,78
2931,78
2932,78
2933,78
2934,78
2935,78
2936,78
2937,78
2938,78
2939,78
2940,78
2941,78
2942,78
2943,78
2944,78
2945,78
2946,78
2947,78
2948,78
2949,78
2950,78
2951,78
2952,78
2953,78
2954,78
2955,78
2956,79
2957,79
2958,79
2959,79
2960,79
2961,79
2962,79
2963,79
2964,79
2965,79
2966,79
2967,79
2968,79
2969,79
2970,79
2971,79
2972,79
2973,79
2974,79
2975,79
2976,79
2977,79
2978,79
2979,79
2980,79
2981,79
2982,79
2983,79
2984,79
2985,79
2986,79
2987,79
2988,79
2989,79
2990,79
2991,79
