0,0
1,0
2,0
3,0
4,0
5,0
6,0
7,0
8,0
9,0
10,0
11,0
12,0
13,0
14,0
15,0
16,0
17,0
18,0
19,0
20,0
21,0
22,0
23,0
24,0
25,0
26,0
27,0
28,0
29,0
30,0
31,0
32,0
33,0
34,0
35,0
36,0
37,0
38,1
39,1
40,1
41,1
42,1
43,1
44,1
45,1
46,1
47,1
48,1
49,1
50,1
51,1
52,1
53,1
54,1
55,1
56,1
57,1
58,1
59,1
60,1
61,1
62,1
63,1
64,1
65,1
66,1
67,1
68,1
69,1
70,1
71,1
72,1
73,1
74,1
75,1
76,2
77,2
78,2
79,2
80,2
81,2
82,2
83,2
84,2
85,2
86,2
87,2
88,2
89,2
90,2
91,2
92,2
93,2
94,2
95,2
96,2
97,2
98,2
99,2
100,2
101,2
102,2
103,2
104,2
105,2
106,2
107,2
108,2
109,2
110,2
111,2
112,2
113,2
114,3
115,3
116,3
117,3
118,3
119,3
120,3
121,3
122,3
123,3
124,3
125,3
126,3
127,3
128,3
129,3
130,3
131,3
132,3
133,3
134,3
135,3
136,3
137,3
138,3
139,3
140,3
141,3
142,3
143,3
144,3
145,3
146,3
147,3
148,3
149,3
150,3
151,3
152,4
153,4
154,4
155,4
156,4
157,4
158,4
159,4
160,4
161,4
162,4
163,4
164,4
165,4
166,4
167,4
168,4
169,4
170,4
171,4
172,4
173,4
174,4
175,4
176,4
177,4
178,4
179,4
180,4
181,4
182,4
183,4
184,4
185,4
186,4
187,4
188,4
189,4
190,5
191,5
192,5
193,5
194,5
195,5
196,5
197,5
198,5
199,5
200,5
201,5
202,5
203,5
204,5
205,5
206,5
207,5
208,5
209,5
210,5
211,5
212,5
213,5
214,5
215,5
216,5
217,5
218,5
219,5
220,5
221,5
222,5
223,5
224,5
225,5
226,5
227,5
228,6
229,6
230,6
231,6
232,6
233,6
234,6
235,6
236,6
237,6
238,6
239,6
240,6
241,6
242,6
243,6
244,6
245,6
246,6
247,6
248,6
249,6
250,6
251,6
252,6
253,6
254,6
255,6
256,6
257,6
258,6
259,6
260,6
261,6
262,6
263,6
264,6
265,6
266,7
267,7
268,7
269,7
270,7
271,7
272,7
273,7
274,7
275,7
276,7
277,7
278,7
279,7
280,7
281,7
282,7
283,7
284,7
285,7
286,7
287,7
288,7
289,7
290,7
291,7
292,7
293,7
294,7
295,7
296,7
297,7
298,7
299,7
300,7
301,7
302,7
303,7
304,8
305,8
306,8
307,8
308,8
309,8
310,8
311,8
312,8
313,8
314,8
315,8
316,8
317,8
318,8
319,8
320,8
321,8
322,8
323,8
324,8
325,8
326,8
327,8
328,8
329,8
330,8
331,8
332,8
333,8
334,8
335,8
336,8
337,8
338,8
339,8
340,8
341,8
342,9
343,9
344,9
345,9
346,9
347,9
348,9
349,9
350,9
351,9
352,9
353,9
354,9
355,9
356,9
357,9
358,9
359,9
360,9
361,9
362,9
363,9
364,9
365,9
366,9
367,9
368,9
369,9
370,9
371,9
372,9
373,9
374,9
375,9
376,9
377,9
378,9
379,9
380,10
381,10
382,10
383,10
384,10
385,10
386,10
387,10
388,10
389,10
390,10
391,10
392,10
393,10
394,10
395,10
396,10
397,10
398,10
399,10
400,10
401,10
402,10
403,10
404,10
405,10
406,10
407,10
408,10
409,10
410,10
411,10
412,10
413,10
414,10
415,10
416,10
417,10
418,11
419,11
420,11
421,11
422,11
423,11
424,11
425,11
426,11
427,11
428,11
429,11
430,11
431,11
432,11
433,11
434,11
435,11
436,11
437,11
438,11
439,11
440,11
441,11
442,11
443,11
444,11
445,11
446,11
447,11
448,11
449,11
450,11
451,11
452,11
453,11
454,11
455,11
456,12
457,12
458,12
459,12
460,12
461,12
462,12
463,12
464,12
465,12
466,12
467,12
468,12
469,12
470,12
471,12
472,12
473,12
474,12
475,12
476,12
477,12
478,12
479,12
480,12
481,12
482,12
483,12
484,12
485,12
486,12
487,12
488,12
489,12
490,12
491,12
492,12
493,12
494,13
495,13
496,13
497,13
498,13
499,13
500,13
501,13
502,13
503,13
504,13
505,13
506,13
507,13
508,13
509,13
510,13
511,13
512,13
513,13
514,13
515,13
516,13
517,13
518,13
519,13
520,13
521,13
522,13
523,13
524,13
525,13
526,13
527,13
528,13
529,13
530,13
531,13
532,14
533,14
534,14
535,14
536,14
537,14
538,14
539,14
540,14
541,14
542,14
543,14
544,14
545,14
546,14
547,14
548,14
549,14
550,14
551,14
552,14
553,14
554,14
555,14
556,14
557,14
558,14
559,14
560,14
561,14
562,14
563,14
564,14
565,14
566,14
567,14
568,14
569,14
570,15
571,15
572,15
573,15
574,15
575,15
576,15
577,15
578,15
579,15
580,15
581,15
582,15
583,15
584,15
585,15
586,15
587,15
588,15
589,15
590,15
591,15
592,15
593,15
594,15
595,15
596,15
597,15
598,15
599,15
600,15
601,15
602,15
603,15
604,15
605,15
606,15
607,15
608,16
609,16
610,16
611,16
612,16
613,16
614,16
615,16
616,16
617,16
618,16
619,16
620,16
621,16
622,16
623,16
624,16
625,16
626,16
627,16
628,16
629,16
630,16
631,16
632,16
633,16
634,16
635,16
636,16
637,16
638,16
639,16
640,16
641,16
642,16
643,16
644,16
645,16
646,17
647,17
648,17
649,17
650,17
651,17
652,17
653,17
654,17
655,17
656,17
657,17
658,17
659,17
660,17
661,17
662,17
663,17
664,17
665,17
666,17
667,17
668,17
669,17
670,17
671,17
672,17
673,17
674,17
675,17
676,17
677,17
678,17
679,17
680,17
681,17
682,17
683,17
684,18
685,18
686,18
687,18
688,18
689,18
690,18
691,18
692,18
693,18
694,18
695,18
696,18
697,18
698,18
699,18
700,18
701,18
702,18
703,18
704,18
705,18
706,18
707,18
708,18
709,18
710,18
711,18
712,18
713,18
714,18
715,18
716,18
717,18
718,18
719,18
720,18
721,18
722,19
723,19
724,19
725,19
726,19
727,19
728,19
729,19
730,19
731,19
732,19
733,19
734,19
735,19
736,19
737,19
738,19
739,19
740,19
741,19
742,19
743,19
744,19
745,19
746,19
747,19
748,19
749,19
750,19
751,19
752,19
753,19
754,19
755,19
756,19
757,19
758,19
759,19
760,20
761,20
762,20
763,20
764,20
765,20
766,20
767,20
768,20
769,20
770,20
771,20
772,20
773,20
774,20
775,20
776,20
777,20
778,20
779,20
780,20
781,20
782,20
783,20
784,20
785,20
786,20
787,20
788,20
789,20
790,20
791,20
792,20
793,20
794,20
795,20
796,20
797,20
798,21
799,21
800,21
801,21
802,21
803,21
804,21
805,21
806,21
807,21
808,21
809,21
810,21
811,21
812,21
813,21
814,21
815,21
816,21
817,21
818,21
819,21
820,21
821,21
822,21
823,21
824,21
825,21
826,21
827,21
828,21
829,21
830,21
831,21
832,21
833,21
834,21
835,21
836,22
837,22
838,22
839,22
840,22
841,22
842,22
843,22
844,22
845,22
846,22
847,22
848,22
849,22
850,22
851,22
852,22
853,22
854,22
855,22
856,22
857,22
858,22
859,22
860,22
861,22
862,22
863,22
864,22
865,22
866,22
867,22
868,22
869,22
870,22
871,22
872,22
873,22
874,23
875,23
876,23
877,23
878,23
879,23
880,23
881,23
882,23
883,23
884,23
885,23
886,23
887,23
888,23
889,23
890,23
891,23
892,23
893,23
894,23
895,23
896,23
897,23
898,23
899,23
900,23
901,23
902,23
903,23
904,23
905,23
906,23
907,23
908,23
909,23
910,23
911,23
912,24
913,24
914,24
915,24
916,24
917,24
918,24
919,24
920,24
921,24
922,24
923,24
924,24
925,24
926,24
927,24
928,24
929,24
930,24
931,24
932,24
933,24
934,24
935,24
936,24
937,24
938,24
939,24
940,24
941,24
942,24
943,24
944,24
945,24
946,24
947,24
948,24
949,24
950,25
951,25
952,25
953,25
954,25
955,25
956,25
957,25
958,25
959,25
960,25
961,25
962,25
963,25
964,25
965,25
966,25
967,25
968,25
969,25
970,25
971,25
972,25
973,25
974,25
975,25
976,25
977,25
978,25
979,25
980,25
981,25
982,25
983,25
984,25
985,25
986,25
987,25
988,26
989,26
990,26
991,26
992,26
993,26
994,26
995,26
996,26
997,26
998,26
999,26
1000,26
1001,26
1002,26
1003,26
1004,26
1005,26
1006,26
1007,26
1008,26
1009,26
1010,26
1011,26
1012,26
1013,26
1014,26
1015,26
1016,26
1017,26
1018,26
1019,26
1020,26
1021,26
1022,26
1023,26
1024,26
1025,26
1026,27
1027,27
1028,27
1029,27
1030,27
1031,27
1032,27
1033,27
1034,27
1035,27
1036,27
1037,27
1038,27
1039,27
1040,27
1041,27
1042,27
1043,27
1044,27
1045,27
1046,27
1047,27
1048,27
1049,27
1050,27
1051,27
1052,27
1053,27
1054,27
1055,27
1056,27
1057,27
1058,27
1059,27
1060,27
1061,27
1062,27
1063,27
1064,28
1065,28
1066,28
1067,28
1068,28
1069,28
1070,28
1071,28
1072,28
1073,28
1074,28
1075,28
1076,28
1077,28
1078,28
1079,28
1080,28
1081,28
1082,28
1083,28
1084,28
1085,28
1086,28
1087,28
1088,28
1089,28
1090,28
1091,28
1092,28
1093,28
1094,28
1095,28
1096,28
1097,28
1098,28
1099,28
1100,28
1101,28
1102,29
1103,29
1104,29
1105,29
1106,29
1107,29
1108,29
1109,29
1110,29
1111,29
1112,29
1113,29
1114,29
1115,29
1116,29
1117,29
1118,29
1119,29
1120,29
1121,29
1122,29
1123,29
1124,29
1125,29
1126,29
1127,29
1128,29
1129,29
1130,29
1131,29
1132,29
1133,29
1134,29
1135,29
1136,29
1137,29
1138,29
1139,29
1140,30
1141,30
1142,30
1143,30
1144,30
1145,30
1146,30
1147,30
1148,30
1149,30
1150,30
1151,30
1152,30
1153,30
1154,30
1155,30
1156,30
1157,30
1158,30
1159,30
1160,30
1161,30
1162,30
1163,30
1164,30
1165,30
1166,30
1167,30
1168,30
1169,30
1170,30
1171,30
1172,30
1173,30
1174,30
1175,30
1176,30
1177,30
1178,31
1179,31
1180,31
1181,31
1182,31
1183,31
1184,31
1185,31
1186,31
1187,31
1188,31
1189,31
1190,31
1191,31
1192,31
1193,31
1194,31
1195,31
1196,31
1197,31
1198,31
1199,31
1200,31
1201,31
1202,31
1203,31
1204,31
1205,31
1206,31
1207,31
1208,31
1209,31
1210,31
1211,31
1212,31
1213,31
1214,31
1215,31
1216,32
1217,32
1218,32
1219,32
1220,32
1221,32
1222,32
1223,32
1224,32
1225,32
1226,32
1227,32
1228,32
1229,32
1230,32
1231,32
1232,32
1233,32
1234,32
1235,32
1236,32
1237,32
1238,32
1239,32
1240,32
1241,32
1242,32
1243,32
1244,32
1245,32
1246,32
1247,32
1248,32
1249,32
1250,32
1251,32
1252,32
1253,32
1254,33
1255,33
1256,33
1257,33
1258,33
1259,33
1260,33
1261,33
1262,33
1263,33
1264,33
1265,33
1266,33
1267,33
1268,33
1269,33
1270,33
1271,33
1272,33
1273,33
1274,33
1275,33
1276,33
1277,33
1278,33
1279,33
1280,33
1281,33
1282,33
1283,33
1284,33
1285,33
1286,33
1287,33
1288,33
1289,33
1290,33
1291,33
1292,34
1293,34
1294,34
1295,34
1296,34
1297,34
1298,34
1299,34
1300,34
1301,34
1302,34
1303,34
1304,34
1305,34
1306,34
1307,34
1308,34
1309,34
1310,34
1311,34
1312,34
1313,34
1314,34
1315,34
1316,34
1317,34
1318,34
1319,34
1320,34
1321,34
1322,34
1323,34
1324,34
1325,34
1326,34
1327,34
1328,34
1329,34
1330,35
1331,35
1332,35
1333,35
1334,35
1335,35
1336,35
1337,35
1338,35
1339,35
1340,35
1341,35
1342,35
1343,35
1344,35
1345,35
1346,35
1347,35
1348,35
1349,35
1350,35
1351,35
1352,35
1353,35
1354,35
1355,35
1356,35
1357,35
1358,35
1359,35
1360,35
1361,35
1362,35
1363,35
1364,35
1365,35
1366,35
1367,35
1368,36
1369,36
1370,36
1371,36
1372,36
1373,36
1374,36
1375,36
1376,36
1377,36
1378,36
1379,36
1380,36
1381,36
1382,36
1383,36
1384,36
1385,36
1386,36
1387,36
1388,36
1389,36
1390,36
1391,36
1392,36
1393,36
1394,36
1395,36
1396,36
1397,36
1398,36
1399,36
1400,36
1401,36
1402,36
1403,36
1404,36
1405,36
1406,37
1407,37
1408,37
1409,37
1410,37
1411,37
1412,37
1413,37
1414,37
1415,37
1416,37
1417,37
1418,37
1419,37
1420,37
1421,37
1422,37
1423,37
1424,37
1425,37
1426,37
1427,37
1428,37
1429,37
1430,37
1431,37
1432,37
1433,37
1434,37
1435,37
1436,37
1437,37
1438,37
1439,37
1440,37
1441,37
1442,37
1443,37
1444,38
1445,38
1446,38
1447,38
1448,38
1449,38
1450,38
1451,38
1452,38
1453,38
1454,38
1455,38
1456,38
1457,38
1458,38
1459,38
1460,38
1461,38
1462,38
1463,38
1464,38
1465,38
1466,38
1467,38
1468,38
1469,38
1470,38
1471,38
1472,38
1473,38
1474,38
1475,38
1476,38
1477,38
1478,38
1479,38
1480,38
1481,38
1482,39
1483,39
1484,39
1485,39
1486,39
1487,39
1488,39
1489,39
1490,39
1491,39
1492,39
1493,39
1494,39
1495,39
1496,39
1497,39
1498,39
1499,39
1500,39
1501,39
1502,39
1503,39
1504,39
1505,39
1506,39
1507,39
1508,39
1509,39
1510,39
1511,39
1512,39
1513,39
1514,39
1515,39
1516,39
1517,39
1518,39
1519,39
1520,40
1521,40
1522,40
1523,40
1524,40
1525,40
1526,40
1527,40
1528,40
1529,40
1530,40
1531,40
1532,40
1533,40
1534,40
1535,40
1536,40
1537,40
1538,40
1539,40
1540,40
1541,40
1542,40
1543,40
1544,40
1545,40
1546,40
1547,40
1548,40
1549,40
1550,40
1551,40
1552,40
1553,40
1554,40
1555,40
1556,40
1557,40
1558,41
1559,41
1560,41
1561,41
1562,41
1563,41
1564,41
1565,41
1566,41
1567,41
1568,41
1569,41
1570,41
1571,41
1572,41
1573,41
1574,41
1575,41
1576,41
1577,41
1578,41
1579,41
1580,41
1581,41
1582,41
1583,41
1584,41
1585,41
1586,41
1587,41
1588,41
1589,41
1590,41
1591,41
1592,41
1593,41
1594,41
1595,41
1596,42
1597,42
1598,42
1599,42
1600,42
1601,42
1602,42
1603,42
1604,42
1605,42
1606,42
1607,42
1608,42
1609,42
1610,42
1611,42
1612,42
1613,42
1614,42
1615,42
1616,42
1617,42
1618,42
1619,42
1620,42
1621,42
1622,42
1623,42
1624,42
1625,42
1626,42
1627,42
1628,42
1629,42
1630,42
1631,42
1632,42
1633,42
1634,43
1635,43
1636,43
1637,43
1638,43
1639,43
1640,43
1641,43
1642,43
1643,43
1644,43
1645,43
1646,43
1647,43
1648,43
1649,43
1650,43
1651,43
1652,43
1653,43
1654,43
1655,43
1656,43
1657,43
1658,43
1659,43
1660,43
1661,43
1662,43
1663,43
1664,43
1665,43
1666,43
1667,43
1668,43
1669,43
1670,43
1671,43
1672,44
1673,44
1674,44
1675,44
1676,44
1677,44
1678,44
1679,44
1680,44
1681,44
1682,44
1683,44
1684,44
1685,44
1686,44
1687,44
1688,44
1689,44
1690,44
1691,44
1692,44
1693,44
1694,44
1695,44
1696,44
1697,44
1698,44
1699,44
1700,44
1701,44
1702,44
1703,44
1704,44
1705,44
1706,44
1707,44
1708,44
1709,44
1710,45
1711,45
1712,45
1713,45
1714,45
1715,45
1716,45
1717,45
1718,45
1719,45
1720,45
1721,45
1722,45
1723,45
1724,45
1725,45
1726,45
1727,45
1728,45
1729,45
1730,45
1731,45
1732,45
1733,45
1734,45
1735,45
1736,45
1737,45
1738,45
1739,45
1740,45
1741,45
1742,45
1743,45
1744,45
1745,45
1746,45
1747,45
1748,46
1749,46
1750,46
1751,46
1752,46
1753,46
1754,46
1755,46
1756,46
1757,46
1758,46
1759,46
1760,46
1761,46
1762,46
1763,46
1764,46
1765,46
1766,46
1767,46
1768,46
1769,46
1770,46
1771,46
1772,46
1773,46
1774,46
1775,46
1776,46
1777,46
1778,46
1779,46
1780,46
1781,46
1782,46
1783,46
1784,46
1785,46
1786,47
1787,47
1788,47
1789,47
1790,47
1791,47
1792,47
1793,47
1794,47
1795,47
1796,47
1797,47
1798,47
1799,47
1800,47
1801,47
1802,47
1803,47
1804,47
1805,47
1806,47
1807,47
1808,47
1809,47
1810,47
1811,47
1812,47
1813,47
1814,47
1815,47
1816,47
1817,47
1818,47
1819,47
1820,47
1821,47
1822,47
1823,47
1824,48
1825,48
1826,48
1827,48
1828,48
1829,48
1830,48
1831,48
1832,48
1833,48
1834,48
1835,48
1836,48
1837,48
1838,48
1839,48
1840,48
1841,48
1842,48
1843,48
1844,48
1845,48
1846,48
1847,48
1848,48
1849,48
1850,48
1851,48
1852,48
1853,48
1854,48
1855,48
1856,48
1857,48
1858,48
1859,48
1860,48
1861,48
1862,48
1863,49
1864,49
1865,49
1866,49
1867,49
1868,49
1869,49
1870,49
1871,49
1872,49
1873,49
1874,49
1875,49
1876,49
1877,49
1878,49
1879,49
1880,49
1881,49
1882,49
1883,49
1884,49
1885,49
1886,49
1887,49
1888,49
1889,49
1890,49
1891,49
1892,49
1893,49
1894,49
1895,49
1896,49
1897,49
1898,49
1899,49
1900,49
1901,49
1902,50
1903,50
1904,50
1905,50
1906,50
1907,50
1908,50
1909,50
1910,50
1911,50
1912,50
1913,50
1914,50
1915,50
1916,50
1917,50
1918,50
1919,50
1920,50
1921,50
1922,50
1923,50
1924,50
1925,50
1926,50
1927,50
1928,50
1929,50
1930,50
1931,50
1932,50
1933,50
1934,50
1935,50
1936,50
1937,50
1938,50
1939,50
1940,50
1941,51
1942,51
1943,51
1944,51
1945,51
1946,51
1947,51
1948,51
1949,51
1950,51
1951,51
1952,51
1953,51
1954,51
1955,51
1956,51
1957,51
1958,51
1959,51
1960,51
1961,51
1962,51
1963,51
1964,51
1965,51
1966,51
1967,51
1968,51
1969,51
1970,51
1971,51
1972,51
1973,51
1974,51
1975,51
1976,51
1977,51
1978,51
1979,51
1980,52
1981,52
1982,52
1983,52
1984,52
1985,52
1986,52
1987,52
1988,52
1989,52
1990,52
1991,52
1992,52
1993,52
1994,52
1995,52
1996,52
1997,52
1998,52
1999,52
2000,52
2001,52
2002,52
2003,52
2004,52
2005,52
2006,52
2007,52
2008,52
2009,52
2010,52
2011,52
2012,52
2013,52
2014,52
2015,52
2016,52
2017,52
2018,52
2019,53
2020,53
2021,53
2022,53
2023,53
2024,53
2025,53
2026,53
2027,53
2028,53
2029,53
2030,53
2031,53
2032,53
2033,53
2034,53
2035,53
2036,53
2037,53
2038,53
2039,53
2040,53
2041,53
2042,53
2043,53
2044,53
2045,53
2046,53
2047,53
2048,53
2049,53
2050,53
2051,53
2052,53
2053,53
2054,53
2055,53
2056,53
2057,53
2058,54
2059,54
2060,54
2061,54
2062,54
2063,54
2064,54
2065,54
2066,54
2067,54
2068,54
2069,54
2070,54
2071,54
2072,54
2073,54
2074,54
2075,54
2076,54
2077,54
2078,54
2079,54
2080,54
2081,54
2082,54
2083,54
2084,54
2085,54
2086,54
2087,54
2088,54
2089,54
2090,54
2091,54
2092,54
2093,54
2094,54
2095,54
2096,54
2097,55
2098,55
2099,55
2100,55
2101,55
2102,55
2103,55
2104,55
2105,55
2106,55
2107,55
2108,55
2109,55
2110,55
2111,55
2112,55
2113,55
2114,55
2115,55
2116,55
2117,55
2118,55
2119,55
2120,55
2121,55
2122,55
2123,55
2124,55
2125,55
2126,55
2127,55
2128,55
2129,55
2130,55
2131,55
2132,55
2133,55
2134,55
2135,55
2136,56
2137,56
2138,56
2139,56
2140,56
2141,56
2142,56
2143,56
2144,56
2145,56
2146,56
2147,56
2148,56
2149,56
2150,56
2151,56
2152,56
2153,56
2154,56
2155,56
2156,56
2157,56
2158,56
2159,56
2160,56
2161,56
2162,56
2163,56
2164,56
2165,56
2166,56
2167,56
2168,56
2169,56
2170,56
2171,56
2172,56
2173,56
2174,56
2175,57
2176,57
2177,57
2178,57
2179,57
2180,57
2181,57
2182,57
2183,57
2184,57
2185,57
2186,57
2187,57
2188,57
2189,57
2190,57
2191,57
2192,57
2193,57
2194,57
2195,57
2196,57
2197,57
2198,57
2199,57
2200,57
2201,57
2202,57
2203,57
2204,57
2205,57
2206,57
2207,57
2208,57
2209,57
2210,57
2211,57
2212,57
2213,57
2214,58
2215,58
2216,58
2217,58
2218,58
2219,58
2220,58
2221,58
2222,58
2223,58
2224,58
2225,58
2226,58
2227,58
2228,58
2229,58
2230,58
2231,58
2232,58
2233,58
2234,58
2235,58
2236,58
2237,58
2238,58
2239,58
2240,58
2241,58
2242,58
2243,58
2244,58
2245,58
2246,58
2247,58
2248,58
2249,58
2250,58
2251,58
2252,58
2253,59
2254,59
2255,59
2256,59
2257,59
2258,59
2259,59
2260,59
2261,59
2262,59
2263,59
2264,59
2265,59
2266,59
2267,59
2268,59
2269,59
2270,59
2271,59
2272,59
2273,59
2274,59
2275,59
2276,59
2277,59
2278,59
2279,59
2280,59
2281,59
2282,59
2283,59
2284,59
2285,59
2286,59
2287,59
2288,59
2289,59
2290,59
2291,59
2292,60
2293,60
2294,60
2295,60
2296,60
2297,60
2298,60
2299,60
2300,60
2301,60
2302,60
2303,60
2304,60
2305,60
2306,60
2307,60
2308,60
2309,60
2310,60
2311,60
2312,60
2313,60
2314,60
2315,60
2316,60
2317,60
2318,60
2319,60
2320,60
2321,60
2322,60
2323,60
2324,60
2325,60
2326,60
2327,60
2328,60
2329,60
2330,60
2331,61
2332,61
2333,61
2334,61
2335,61
2336,61
2337,61
2338,61
2339,61
2340,61
2341,61
2342,61
2343,61
2344,61
2345,61
2346,61
2347,61
2348,61
2349,61
2350,61
2351,61
2352,61
2353,61
2354,61
2355,61
2356,61
2357,61
2358,61
2359,61
2360,61
2361,61
2362,61
2363,61
2364,61
2365,61
2366,61
2367,61
2368,61
2369,61
2370,62
2371,62
2372,62
2373,62
2374,62
2375,62
2376,62
2377,62
2378,62
2379,62
2380,62
2381,62
2382,62
2383,62
2384,62
2385,62
2386,62
2387,62
2388,62
2389,62
2390,62
2391,62
2392,62
2393,62
2394,62
2395,62
2396,62
2397,62
2398,62
2399,62
2400,62
2401,62
2402,62
2403,62
2404,62
2405,62
2406,62
2407,62
2408,62
2409,63
2410,63
2411,63
2412,63
2413,63
2414,63
2415,63
2416,63
2417,63
2418,63
2419,63
2420,63
2421,63
2422,63
2423,63
2424,63
2425,63
2426,63
2427,63
2428,63
2429,63
2430,63
2431,63
2432,63
2433,63
2434,63
2435,63
2436,63
2437,63
2438,63
2439,63
2440,63
2441,63
2442,63
2443,63
2444,63
2445,63
2446,63
2447,63
2448,64
2449,64
2450,64
2451,64
2452,64
2453,64
2454,64
2455,64
2456,64
2457,64
2458,64
2459,64
2460,64
2461,64
2462,64
2463,64
2464,64
2465,64
2466,64
2467,64
2468,64
2469,64
2470,64
2471,64
2472,64
2473,64
2474,64
2475,64
2476,64
2477,64
2478,64
2479,64
2480,64
2481,64
2482,64
2483,64
2484,64
2485,64
2486,64
2487,65
2488,65
2489,65
2490,65
2491,65
2492,65
2493,65
2494,65
2495,65
2496,65
2497,65
2498,65
2499,65
2500,65
2501,65
2502,65
2503,65
2504,65
2505,65
2506,65
2507,65
2508,65
2509,65
2510,65
2511,65
2512,65
2513,65
2514,65
2515,65
2516,65
2517,65
2518,65
2519,65
2520,65
2521,65
2522,65
2523,65
2524,65
2525,65
2526,66
2527,66
2528,66
2529,66
2530,66
2531,66
2532,66
2533,66
2534,66
2535,66
2536,66
2537,66
2538,66
2539,66
2540,66
2541,66
2542,66
2543,66
2544,66
2545,66
2546,66
2547,66
2548,66
2549,66
2550,66
2551,66
2552,66
2553,66
2554,66
2555,66
2556,66
2557,66
2558,66
2559,66
2560,66
2561,66
2562,66
2563,66
2564,66
2565,67
2566,67
2567,67
2568,67
2569,67
2570,67
2571,67
2572,67
2573,67
2574,67
2575,67
2576,67
2577,67
2578,67
2579,67
2580,67
2581,67
2582,67
2583,67
2584,67
2585,67
2586,67
2587,67
2588,67
2589,67
2590,67
2591,67
2592,67
2593,67
2594,67
2595,67
2596,67
2597,67
2598,67
2599,67
2600,67
2601,67
2602,67
2603,67
2604,68
2605,68
2606,68
2607,68
2608,68
2609,68
2610,68
2611,68
2612,68
2613,68
2614,68
2615,68
2616,68
2617,68
2618,68
2619,68
2620,68
2621,68
2622,68
2623,68
2624,68
2625,68
2626,68
2627,68
2628,68
2629,68
2630,68
2631,68
2632,68
2633,68
2634,68
2635,68
2636,68
2637,68
2638,68
2639,68
2640,68
2641,68
2642,68
2643,69
2644,69
2645,69
2646,69
2647,69
2648,69
2649,69
2650,69
2651,69
2652,69
2653,69
2654,69
2655,69
2656,69
2657,69
2658,69
2659,69
2660,69
2661,69
2662,69
2663,69
2664,69
2665,69
2666,69
2667,69
2668,69
2669,69
2670,69
2671,69
2672,69
2673,69
2674,69
2675,69
2676,69
2677,69
2678,69
2679,69
2680,69
2681,69
2682,70
2683,70
2684,70
2685,70
2686,70
2687,70
2688,70
2689,70
2690,70
2691,70
2692,70
2693,70
2694,70
2695,70
2696,70
2697,70
2698,70
2699,70
2700,70
2701,70
2702,70
2703,70
2704,70
2705,70
2706,70
2707,70
2708,70
2709,70
2710,70
2711,70
2712,70
2713,70
2714,70
2715,70
2716,70
2717,70
2718,70
2719,70
2720,70
2721,71
2722,71
2723,71
2724,71
2725,71
2726,71
2727,71
2728,71
2729,71
2730,71
2731,71
2732,71
2733,71
2734,71
2735,71
2736,71
2737,71
2738,71
2739,71
2740,71
2741,71
2742,71
2743,71
2744,71
2745,71
2746,71
2747,71
2748,71
2749,71
2750,71
2751,71
2752,71
2753,71
2754,71
2755,71
2756,71
2757,71
2758,71
2759,71
2760,72
2761,72
2762,72
2763,72
2764,72
2765,72
2766,72
2767,72
2768,72
2769,72
2770,72
2771,72
2772,72
2773,72
2774,72
2775,72
2776,72
2777,72
2778,72
2779,72
2780,72
2781,72
2782,72
2783,72
2784,72
2785,72
2786,72
2787,72
2788,72
2789,72
2790,72
2791,72
2792,72
2793,72
2794,72
2795,72
2796,72
2797,72
2798,72
2799,73
2800,73
2801,73
2802,73
2803,73
2804,73
2805,73
2806,73
2807,73
2808,73
2809,73
2810,73
2811,73
2812,73
2813,73
2814,73
2815,73
2816,73
2817,73
2818,73
2819,73
2820,73
2821,73
2822,73
2823,73
2824,73
2825,73
2826,73
2827,73
2828,73
2829,73
2830,73
2831,73
2832,73
2833,73
2834,73
2835,73
2836,73
2837,73
2838,74
2839,74
2840,74
2841,74
2842,74
2843,74
2844,74
2845,74
2846,74
2847,74
2848,74
2849,74
2850,74
2851,74
2852,74
2853,74
2854,74
2855,74
2856,74
2857,74
2858,74
2859,74
2860,74
2861,74
2862,74
2863,74
2864,74
2865,74
2866,74
2867,74
2868,74
2869,74
2870,74
2871,74
2872,74
2873,74
2874,74
2875,74
2876,74
2877,75
2878,75
2879,75
2880,75
2881,75
2882,75
2883,75
2884,75
2885,75
2886,75
2887,75
2888,75
2889,75
2890,75
2891,75
2892,75
2893,75
2894,75
2895,75
2896,75
2897,75
2898,75
2899,75
2900,75
2901,75
2902,75
2903,75
2904,75
2905,75
2906,75
2907,75
2908,75
2909,75
2910,75
2911,75
2912,75
2913,75
2914,75
2915,75
2916,76
2917,76
2918,76
2919,76
2920,76
2921,76
2922,76
2923,76
2924,76
2925,76
2926,76
2927,76
2928,76
2929,76
2930,76
2931,76
2932,76
2933,76
2934,76
2935,76
2936,76
2937,76
2938,76
2939,76
2940,76
2941,76
2942,76
2943,76
2944,76
2945,76
2946,76
2947,76
2948,76
2949,76
2950,76
2951,76
2952,76
2953,76
2954,76
2955,77
2956,77
2957,77
2958,77
2959,77
2960,77
2961,77
2962,77
2963,77
2964,77
2965,77
2966,77
2967,77
2968,77
2969,77
2970,77
2971,77
2972,77
2973,77
2974,77
2975,77
2976,77
2977,77
2978,77
2979,77
2980,77
2981,77
2982,77
2983,77
2984,77
2985,77
2986,77
2987,77
2988,77
2989,77
2990,77
2991,77
2992,77
2993,77
2994,78
2995,78
2996,78
2997,78
2998,78
2999,78
3000,78
3001,78
3002,78
3003,78
3004,78
3005,78
3006,78
3007,78
3008,78
3009,78
3010,78
3011,78
3012,78
3013,78
3014,78
3015,78
3016,78
3017,78
3018,78
3019,78
3020,78
3021,78
3022,78
3023,78
3024,78
3025,78
3026,78
3027,78
3028,78
3029,78
3030,78
3031,78
3032,78
3033,79
3034,79
3035,79
3036,79
3037,79
3038,79
3039,79
3040,79
3041,79
3042,79
3043,79
3044,79
3045,79
3046,79
3047,79
3048,79
3049,79
3050,79
3051,79
3052,79
3053,79
3054,79
3055,79
3056,79
3057,79
3058,79
3059,79
3060,79
3061,79
3062,79
3063,79
3064,79
3065,79
3066,79
3067,79
3068,79
3069,79
3070,79
3071,79
