0,0
1,0
2,0
3,0
4,0
5,0
6,0
7,0
8,0
9,0
10,0
11,0
12,0
13,0
14,0
15,0
16,0
17,0
18,0
19,1
20,1
21,1
22,1
23,1
24,1
25,1
26,1
27,1
28,1
29,1
30,1
31,1
32,1
33,1
34,1
35,1
36,1
37,1
38,2
39,2
40,2
41,2
42,2
43,2
44,2
45,2
46,2
47,2
48,2
49,2
50,2
51,2
52,2
53,2
54,2
55,2
56,2
57,3
58,3
59,3
60,3
61,3
62,3
63,3
64,3
65,3
66,3
67,3
68,3
69,3
70,3
71,3
72,3
73,3
74,3
75,3
76,4
77,4
78,4
79,4
80,4
81,4
82,4
83,4
84,4
85,4
86,4
87,4
88,4
89,4
90,4
91,4
92,4
93,4
94,4
95,5
96,5
97,5
98,5
99,5
100,5
101,5
102,5
103,5
104,5
105,5
106,5
107,5
108,5
109,5
110,5
111,5
112,5
113,5
114,6
115,6
116,6
117,6
118,6
119,6
120,6
121,6
122,6
123,6
124,6
125,6
126,6
127,6
128,6
129,6
130,6
131,6
132,6
133,7
134,7
135,7
136,7
137,7
138,7
139,7
140,7
141,7
142,7
143,7
144,7
145,7
146,7
147,7
148,7
149,7
150,7
151,7
152,8
153,8
154,8
155,8
156,8
157,8
158,8
159,8
160,8
161,8
162,8
163,8
164,8
165,8
166,8
167,8
168,8
169,8
170,8
171,9
172,9
173,9
174,9
175,9
176,9
177,9
178,9
179,9
180,9
181,9
182,9
183,9
184,9
185,9
186,9
187,9
188,9
189,9
190,10
191,10
192,10
193,10
194,10
195,10
196,10
197,10
198,10
199,10
200,10
201,10
202,10
203,10
204,10
205,10
206,10
207,10
208,10
209,11
210,11
211,11
212,11
213,11
214,11
215,11
216,11
217,11
218,11
219,11
220,11
221,11
222,11
223,11
224,11
225,11
226,11
227,11
228,12
229,12
230,12
231,12
232,12
233,12
234,12
235,12
236,12
237,12
238,12
239,12
240,12
241,12
242,12
243,12
244,12
245,12
246,12
247,13
248,13
249,13
250,13
251,13
252,13
253,13
254,13
255,13
256,13
257,13
258,13
259,13
260,13
261,13
262,13
263,13
264,13
265,13
266,14
267,14
268,14
269,14
270,14
271,14
272,14
273,14
274,14
275,14
276,14
277,14
278,14
279,14
280,14
281,14
282,14
283,14
284,14
285,15
286,15
287,15
288,15
289,15
290,15
291,15
292,15
293,15
294,15
295,15
296,15
297,15
298,15
299,15
300,15
301,15
302,15
303,15
304,16
305,16
306,16
307,16
308,16
309,16
310,16
311,16
312,16
313,16
314,16
315,16
316,16
317,16
318,16
319,16
320,16
321,16
322,16
323,17
324,17
325,17
326,17
327,17
328,17
329,17
330,17
331,17
332,17
333,17
334,17
335,17
336,17
337,17
338,17
339,17
340,17
341,17
342,18
343,18
344,18
345,18
346,18
347,18
348,18
349,18
350,18
351,18
352,18
353,18
354,18
355,18
356,18
357,18
358,18
359,18
360,18
361,19
362,19
363,19
364,19
365,19
366,19
367,19
368,19
369,19
370,19
371,19
372,19
373,19
374,19
375,19
376,19
377,19
378,19
379,19
380,20
381,20
382,20
383,20
384,20
385,20
386,20
387,20
388,20
389,20
390,20
391,20
392,20
393,20
394,20
395,20
396,20
397,20
398,20
399,21
400,21
401,21
402,21
403,21
404,21
405,21
406,21
407,21
408,21
409,21
410,21
411,21
412,21
413,21
414,21
415,21
416,21
417,21
418,22
419,22
420,22
421,22
422,22
423,22
424,22
425,22
426,22
427,22
428,22
429,22
430,22
431,22
432,22
433,22
434,22
435,22
436,22
437,23
438,23
439,23
440,23
441,23
442,23
443,23
444,23
445,23
446,23
447,23
448,23
449,23
450,23
451,23
452,23
453,23
454,23
455,23
456,24
457,24
458,24
459,24
460,24
461,24
462,24
463,24
464,24
465,24
466,24
467,24
468,24
469,24
470,24
471,24
472,24
473,24
474,24
475,25
476,25
477,25
478,25
479,25
480,25
481,25
482,25
483,25
484,25
485,25
486,25
487,25
488,25
489,25
490,25
491,25
492,25
493,25
494,26
495,26
496,26
497,26
498,26
499,26
500,26
501,26
502,26
503,26
504,26
505,26
506,26
507,26
508,26
509,26
510,26
511,26
512,26
513,27
514,27
515,27
516,27
517,27
518,27
519,27
520,27
521,27
522,27
523,27
524,27
525,27
526,27
527,27
528,27
529,27
530,27
531,27
532,28
533,28
534,28
535,28
536,28
537,28
538,28
539,28
540,28
541,28
542,28
543,28
544,28
545,28
546,28
547,28
548,28
549,28
550,28
551,29
552,29
553,29
554,29
555,29
556,29
557,29
558,29
559,29
560,29
561,29
562,29
563,29
564,29
565,29
566,29
567,29
568,29
569,29
570,30
571,30
572,30
573,30
574,30
575,30
576,30
577,30
578,30
579,30
580,30
581,30
582,30
583,30
584,30
585,30
586,30
587,30
588,30
589,31
590,31
591,31
592,31
593,31
594,31
595,31
596,31
597,31
598,31
599,31
600,31
601,31
602,31
603,31
604,31
605,31
606,31
607,31
608,32
609,32
610,32
611,32
612,32
613,32
614,32
615,32
616,32
617,32
618,32
619,32
620,32
621,32
622,32
623,32
624,32
625,32
626,32
627,32
628,33
629,33
630,33
631,33
632,33
633,33
634,33
635,33
636,33
637,33
638,33
639,33
640,33
641,33
642,33
643,33
644,33
645,33
646,33
647,33
648,34
649,34
650,34
651,34
652,34
653,34
654,34
655,34
656,34
657,34
658,34
659,34
660,34
661,34
662,34
663,34
664,34
665,34
666,34
667,34
668,35
669,35
670,35
671,35
672,35
673,35
674,35
675,35
676,35
677,35
678,35
679,35
680,35
681,35
682,35
683,35
684,35
685,35
686,35
687,35
688,36
689,36
690,36
691,36
692,36
693,36
694,36
695,36
696,36
697,36
698,36
699,36
700,36
701,36
702,36
703,36
704,36
705,36
706,36
707,36
708,37
709,37
710,37
711,37
712,37
713,37
714,37
715,37
716,37
717,37
718,37
719,37
720,37
721,37
722,37
723,37
724,37
725,37
726,37
727,37
728,38
729,38
730,38
731,38
732,38
733,38
734,38
735,38
736,38
737,38
738,38
739,38
740,38
741,38
742,38
743,38
744,38
745,38
746,38
747,38
748,39
749,39
750,39
751,39
752,39
753,39
754,39
755,39
756,39
757,39
758,39
759,39
760,39
761,39
762,39
763,39
764,39
765,39
766,39
767,39
