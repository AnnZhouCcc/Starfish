0,0
1,0
2,0
3,0
4,0
5,0
6,0
7,0
8,0
9,0
10,0
11,0
12,0
13,0
14,0
15,0
16,0
17,0
18,0
19,0
20,0
21,0
22,0
23,0
24,0
25,0
26,0
27,0
28,0
29,0
30,0
31,0
32,0
33,0
34,0
35,0
36,0
37,1
38,1
39,1
40,1
41,1
42,1
43,1
44,1
45,1
46,1
47,1
48,1
49,1
50,1
51,1
52,1
53,1
54,1
55,1
56,1
57,1
58,1
59,1
60,1
61,1
62,1
63,1
64,1
65,1
66,1
67,1
68,1
69,1
70,1
71,1
72,1
73,1
74,2
75,2
76,2
77,2
78,2
79,2
80,2
81,2
82,2
83,2
84,2
85,2
86,2
87,2
88,2
89,2
90,2
91,2
92,2
93,2
94,2
95,2
96,2
97,2
98,2
99,2
100,2
101,2
102,2
103,2
104,2
105,2
106,2
107,2
108,2
109,2
110,2
111,3
112,3
113,3
114,3
115,3
116,3
117,3
118,3
119,3
120,3
121,3
122,3
123,3
124,3
125,3
126,3
127,3
128,3
129,3
130,3
131,3
132,3
133,3
134,3
135,3
136,3
137,3
138,3
139,3
140,3
141,3
142,3
143,3
144,3
145,3
146,3
147,3
148,4
149,4
150,4
151,4
152,4
153,4
154,4
155,4
156,4
157,4
158,4
159,4
160,4
161,4
162,4
163,4
164,4
165,4
166,4
167,4
168,4
169,4
170,4
171,4
172,4
173,4
174,4
175,4
176,4
177,4
178,4
179,4
180,4
181,4
182,4
183,4
184,4
185,5
186,5
187,5
188,5
189,5
190,5
191,5
192,5
193,5
194,5
195,5
196,5
197,5
198,5
199,5
200,5
201,5
202,5
203,5
204,5
205,5
206,5
207,5
208,5
209,5
210,5
211,5
212,5
213,5
214,5
215,5
216,5
217,5
218,5
219,5
220,5
221,5
222,6
223,6
224,6
225,6
226,6
227,6
228,6
229,6
230,6
231,6
232,6
233,6
234,6
235,6
236,6
237,6
238,6
239,6
240,6
241,6
242,6
243,6
244,6
245,6
246,6
247,6
248,6
249,6
250,6
251,6
252,6
253,6
254,6
255,6
256,6
257,6
258,6
259,7
260,7
261,7
262,7
263,7
264,7
265,7
266,7
267,7
268,7
269,7
270,7
271,7
272,7
273,7
274,7
275,7
276,7
277,7
278,7
279,7
280,7
281,7
282,7
283,7
284,7
285,7
286,7
287,7
288,7
289,7
290,7
291,7
292,7
293,7
294,7
295,7
296,8
297,8
298,8
299,8
300,8
301,8
302,8
303,8
304,8
305,8
306,8
307,8
308,8
309,8
310,8
311,8
312,8
313,8
314,8
315,8
316,8
317,8
318,8
319,8
320,8
321,8
322,8
323,8
324,8
325,8
326,8
327,8
328,8
329,8
330,8
331,8
332,8
333,9
334,9
335,9
336,9
337,9
338,9
339,9
340,9
341,9
342,9
343,9
344,9
345,9
346,9
347,9
348,9
349,9
350,9
351,9
352,9
353,9
354,9
355,9
356,9
357,9
358,9
359,9
360,9
361,9
362,9
363,9
364,9
365,9
366,9
367,9
368,9
369,9
370,10
371,10
372,10
373,10
374,10
375,10
376,10
377,10
378,10
379,10
380,10
381,10
382,10
383,10
384,10
385,10
386,10
387,10
388,10
389,10
390,10
391,10
392,10
393,10
394,10
395,10
396,10
397,10
398,10
399,10
400,10
401,10
402,10
403,10
404,10
405,10
406,10
407,11
408,11
409,11
410,11
411,11
412,11
413,11
414,11
415,11
416,11
417,11
418,11
419,11
420,11
421,11
422,11
423,11
424,11
425,11
426,11
427,11
428,11
429,11
430,11
431,11
432,11
433,11
434,11
435,11
436,11
437,11
438,11
439,11
440,11
441,11
442,11
443,11
444,12
445,12
446,12
447,12
448,12
449,12
450,12
451,12
452,12
453,12
454,12
455,12
456,12
457,12
458,12
459,12
460,12
461,12
462,12
463,12
464,12
465,12
466,12
467,12
468,12
469,12
470,12
471,12
472,12
473,12
474,12
475,12
476,12
477,12
478,12
479,12
480,12
481,13
482,13
483,13
484,13
485,13
486,13
487,13
488,13
489,13
490,13
491,13
492,13
493,13
494,13
495,13
496,13
497,13
498,13
499,13
500,13
501,13
502,13
503,13
504,13
505,13
506,13
507,13
508,13
509,13
510,13
511,13
512,13
513,13
514,13
515,13
516,13
517,13
518,14
519,14
520,14
521,14
522,14
523,14
524,14
525,14
526,14
527,14
528,14
529,14
530,14
531,14
532,14
533,14
534,14
535,14
536,14
537,14
538,14
539,14
540,14
541,14
542,14
543,14
544,14
545,14
546,14
547,14
548,14
549,14
550,14
551,14
552,14
553,14
554,14
555,15
556,15
557,15
558,15
559,15
560,15
561,15
562,15
563,15
564,15
565,15
566,15
567,15
568,15
569,15
570,15
571,15
572,15
573,15
574,15
575,15
576,15
577,15
578,15
579,15
580,15
581,15
582,15
583,15
584,15
585,15
586,15
587,15
588,15
589,15
590,15
591,15
592,16
593,16
594,16
595,16
596,16
597,16
598,16
599,16
600,16
601,16
602,16
603,16
604,16
605,16
606,16
607,16
608,16
609,16
610,16
611,16
612,16
613,16
614,16
615,16
616,16
617,16
618,16
619,16
620,16
621,16
622,16
623,16
624,16
625,16
626,16
627,16
628,16
629,17
630,17
631,17
632,17
633,17
634,17
635,17
636,17
637,17
638,17
639,17
640,17
641,17
642,17
643,17
644,17
645,17
646,17
647,17
648,17
649,17
650,17
651,17
652,17
653,17
654,17
655,17
656,17
657,17
658,17
659,17
660,17
661,17
662,17
663,17
664,17
665,17
666,18
667,18
668,18
669,18
670,18
671,18
672,18
673,18
674,18
675,18
676,18
677,18
678,18
679,18
680,18
681,18
682,18
683,18
684,18
685,18
686,18
687,18
688,18
689,18
690,18
691,18
692,18
693,18
694,18
695,18
696,18
697,18
698,18
699,18
700,18
701,18
702,18
703,19
704,19
705,19
706,19
707,19
708,19
709,19
710,19
711,19
712,19
713,19
714,19
715,19
716,19
717,19
718,19
719,19
720,19
721,19
722,19
723,19
724,19
725,19
726,19
727,19
728,19
729,19
730,19
731,19
732,19
733,19
734,19
735,19
736,19
737,19
738,19
739,19
740,20
741,20
742,20
743,20
744,20
745,20
746,20
747,20
748,20
749,20
750,20
751,20
752,20
753,20
754,20
755,20
756,20
757,20
758,20
759,20
760,20
761,20
762,20
763,20
764,20
765,20
766,20
767,20
768,20
769,20
770,20
771,20
772,20
773,20
774,20
775,20
776,20
777,21
778,21
779,21
780,21
781,21
782,21
783,21
784,21
785,21
786,21
787,21
788,21
789,21
790,21
791,21
792,21
793,21
794,21
795,21
796,21
797,21
798,21
799,21
800,21
801,21
802,21
803,21
804,21
805,21
806,21
807,21
808,21
809,21
810,21
811,21
812,21
813,21
814,22
815,22
816,22
817,22
818,22
819,22
820,22
821,22
822,22
823,22
824,22
825,22
826,22
827,22
828,22
829,22
830,22
831,22
832,22
833,22
834,22
835,22
836,22
837,22
838,22
839,22
840,22
841,22
842,22
843,22
844,22
845,22
846,22
847,22
848,22
849,22
850,22
851,23
852,23
853,23
854,23
855,23
856,23
857,23
858,23
859,23
860,23
861,23
862,23
863,23
864,23
865,23
866,23
867,23
868,23
869,23
870,23
871,23
872,23
873,23
874,23
875,23
876,23
877,23
878,23
879,23
880,23
881,23
882,23
883,23
884,23
885,23
886,23
887,23
888,24
889,24
890,24
891,24
892,24
893,24
894,24
895,24
896,24
897,24
898,24
899,24
900,24
901,24
902,24
903,24
904,24
905,24
906,24
907,24
908,24
909,24
910,24
911,24
912,24
913,24
914,24
915,24
916,24
917,24
918,24
919,24
920,24
921,24
922,24
923,24
924,24
925,25
926,25
927,25
928,25
929,25
930,25
931,25
932,25
933,25
934,25
935,25
936,25
937,25
938,25
939,25
940,25
941,25
942,25
943,25
944,25
945,25
946,25
947,25
948,25
949,25
950,25
951,25
952,25
953,25
954,25
955,25
956,25
957,25
958,25
959,25
960,25
961,25
962,26
963,26
964,26
965,26
966,26
967,26
968,26
969,26
970,26
971,26
972,26
973,26
974,26
975,26
976,26
977,26
978,26
979,26
980,26
981,26
982,26
983,26
984,26
985,26
986,26
987,26
988,26
989,26
990,26
991,26
992,26
993,26
994,26
995,26
996,26
997,26
998,26
999,27
1000,27
1001,27
1002,27
1003,27
1004,27
1005,27
1006,27
1007,27
1008,27
1009,27
1010,27
1011,27
1012,27
1013,27
1014,27
1015,27
1016,27
1017,27
1018,27
1019,27
1020,27
1021,27
1022,27
1023,27
1024,27
1025,27
1026,27
1027,27
1028,27
1029,27
1030,27
1031,27
1032,27
1033,27
1034,27
1035,27
1036,28
1037,28
1038,28
1039,28
1040,28
1041,28
1042,28
1043,28
1044,28
1045,28
1046,28
1047,28
1048,28
1049,28
1050,28
1051,28
1052,28
1053,28
1054,28
1055,28
1056,28
1057,28
1058,28
1059,28
1060,28
1061,28
1062,28
1063,28
1064,28
1065,28
1066,28
1067,28
1068,28
1069,28
1070,28
1071,28
1072,28
1073,29
1074,29
1075,29
1076,29
1077,29
1078,29
1079,29
1080,29
1081,29
1082,29
1083,29
1084,29
1085,29
1086,29
1087,29
1088,29
1089,29
1090,29
1091,29
1092,29
1093,29
1094,29
1095,29
1096,29
1097,29
1098,29
1099,29
1100,29
1101,29
1102,29
1103,29
1104,29
1105,29
1106,29
1107,29
1108,29
1109,29
1110,30
1111,30
1112,30
1113,30
1114,30
1115,30
1116,30
1117,30
1118,30
1119,30
1120,30
1121,30
1122,30
1123,30
1124,30
1125,30
1126,30
1127,30
1128,30
1129,30
1130,30
1131,30
1132,30
1133,30
1134,30
1135,30
1136,30
1137,30
1138,30
1139,30
1140,30
1141,30
1142,30
1143,30
1144,30
1145,30
1146,30
1147,31
1148,31
1149,31
1150,31
1151,31
1152,31
1153,31
1154,31
1155,31
1156,31
1157,31
1158,31
1159,31
1160,31
1161,31
1162,31
1163,31
1164,31
1165,31
1166,31
1167,31
1168,31
1169,31
1170,31
1171,31
1172,31
1173,31
1174,31
1175,31
1176,31
1177,31
1178,31
1179,31
1180,31
1181,31
1182,31
1183,31
1184,32
1185,32
1186,32
1187,32
1188,32
1189,32
1190,32
1191,32
1192,32
1193,32
1194,32
1195,32
1196,32
1197,32
1198,32
1199,32
1200,32
1201,32
1202,32
1203,32
1204,32
1205,32
1206,32
1207,32
1208,32
1209,32
1210,32
1211,32
1212,32
1213,32
1214,32
1215,32
1216,32
1217,32
1218,32
1219,32
1220,32
1221,33
1222,33
1223,33
1224,33
1225,33
1226,33
1227,33
1228,33
1229,33
1230,33
1231,33
1232,33
1233,33
1234,33
1235,33
1236,33
1237,33
1238,33
1239,33
1240,33
1241,33
1242,33
1243,33
1244,33
1245,33
1246,33
1247,33
1248,33
1249,33
1250,33
1251,33
1252,33
1253,33
1254,33
1255,33
1256,33
1257,33
1258,34
1259,34
1260,34
1261,34
1262,34
1263,34
1264,34
1265,34
1266,34
1267,34
1268,34
1269,34
1270,34
1271,34
1272,34
1273,34
1274,34
1275,34
1276,34
1277,34
1278,34
1279,34
1280,34
1281,34
1282,34
1283,34
1284,34
1285,34
1286,34
1287,34
1288,34
1289,34
1290,34
1291,34
1292,34
1293,34
1294,34
1295,35
1296,35
1297,35
1298,35
1299,35
1300,35
1301,35
1302,35
1303,35
1304,35
1305,35
1306,35
1307,35
1308,35
1309,35
1310,35
1311,35
1312,35
1313,35
1314,35
1315,35
1316,35
1317,35
1318,35
1319,35
1320,35
1321,35
1322,35
1323,35
1324,35
1325,35
1326,35
1327,35
1328,35
1329,35
1330,35
1331,35
1332,36
1333,36
1334,36
1335,36
1336,36
1337,36
1338,36
1339,36
1340,36
1341,36
1342,36
1343,36
1344,36
1345,36
1346,36
1347,36
1348,36
1349,36
1350,36
1351,36
1352,36
1353,36
1354,36
1355,36
1356,36
1357,36
1358,36
1359,36
1360,36
1361,36
1362,36
1363,36
1364,36
1365,36
1366,36
1367,36
1368,36
1369,37
1370,37
1371,37
1372,37
1373,37
1374,37
1375,37
1376,37
1377,37
1378,37
1379,37
1380,37
1381,37
1382,37
1383,37
1384,37
1385,37
1386,37
1387,37
1388,37
1389,37
1390,37
1391,37
1392,37
1393,37
1394,37
1395,37
1396,37
1397,37
1398,37
1399,37
1400,37
1401,37
1402,37
1403,37
1404,37
1405,37
1406,38
1407,38
1408,38
1409,38
1410,38
1411,38
1412,38
1413,38
1414,38
1415,38
1416,38
1417,38
1418,38
1419,38
1420,38
1421,38
1422,38
1423,38
1424,38
1425,38
1426,38
1427,38
1428,38
1429,38
1430,38
1431,38
1432,38
1433,38
1434,38
1435,38
1436,38
1437,38
1438,38
1439,38
1440,38
1441,38
1442,38
1443,39
1444,39
1445,39
1446,39
1447,39
1448,39
1449,39
1450,39
1451,39
1452,39
1453,39
1454,39
1455,39
1456,39
1457,39
1458,39
1459,39
1460,39
1461,39
1462,39
1463,39
1464,39
1465,39
1466,39
1467,39
1468,39
1469,39
1470,39
1471,39
1472,39
1473,39
1474,39
1475,39
1476,39
1477,39
1478,39
1479,39
1480,40
1481,40
1482,40
1483,40
1484,40
1485,40
1486,40
1487,40
1488,40
1489,40
1490,40
1491,40
1492,40
1493,40
1494,40
1495,40
1496,40
1497,40
1498,40
1499,40
1500,40
1501,40
1502,40
1503,40
1504,40
1505,40
1506,40
1507,40
1508,40
1509,40
1510,40
1511,40
1512,40
1513,40
1514,40
1515,40
1516,40
1517,41
1518,41
1519,41
1520,41
1521,41
1522,41
1523,41
1524,41
1525,41
1526,41
1527,41
1528,41
1529,41
1530,41
1531,41
1532,41
1533,41
1534,41
1535,41
1536,41
1537,41
1538,41
1539,41
1540,41
1541,41
1542,41
1543,41
1544,41
1545,41
1546,41
1547,41
1548,41
1549,41
1550,41
1551,41
1552,41
1553,41
1554,42
1555,42
1556,42
1557,42
1558,42
1559,42
1560,42
1561,42
1562,42
1563,42
1564,42
1565,42
1566,42
1567,42
1568,42
1569,42
1570,42
1571,42
1572,42
1573,42
1574,42
1575,42
1576,42
1577,42
1578,42
1579,42
1580,42
1581,42
1582,42
1583,42
1584,42
1585,42
1586,42
1587,42
1588,42
1589,42
1590,42
1591,43
1592,43
1593,43
1594,43
1595,43
1596,43
1597,43
1598,43
1599,43
1600,43
1601,43
1602,43
1603,43
1604,43
1605,43
1606,43
1607,43
1608,43
1609,43
1610,43
1611,43
1612,43
1613,43
1614,43
1615,43
1616,43
1617,43
1618,43
1619,43
1620,43
1621,43
1622,43
1623,43
1624,43
1625,43
1626,43
1627,43
1628,44
1629,44
1630,44
1631,44
1632,44
1633,44
1634,44
1635,44
1636,44
1637,44
1638,44
1639,44
1640,44
1641,44
1642,44
1643,44
1644,44
1645,44
1646,44
1647,44
1648,44
1649,44
1650,44
1651,44
1652,44
1653,44
1654,44
1655,44
1656,44
1657,44
1658,44
1659,44
1660,44
1661,44
1662,44
1663,44
1664,44
1665,45
1666,45
1667,45
1668,45
1669,45
1670,45
1671,45
1672,45
1673,45
1674,45
1675,45
1676,45
1677,45
1678,45
1679,45
1680,45
1681,45
1682,45
1683,45
1684,45
1685,45
1686,45
1687,45
1688,45
1689,45
1690,45
1691,45
1692,45
1693,45
1694,45
1695,45
1696,45
1697,45
1698,45
1699,45
1700,45
1701,45
1702,46
1703,46
1704,46
1705,46
1706,46
1707,46
1708,46
1709,46
1710,46
1711,46
1712,46
1713,46
1714,46
1715,46
1716,46
1717,46
1718,46
1719,46
1720,46
1721,46
1722,46
1723,46
1724,46
1725,46
1726,46
1727,46
1728,46
1729,46
1730,46
1731,46
1732,46
1733,46
1734,46
1735,46
1736,46
1737,46
1738,46
1739,47
1740,47
1741,47
1742,47
1743,47
1744,47
1745,47
1746,47
1747,47
1748,47
1749,47
1750,47
1751,47
1752,47
1753,47
1754,47
1755,47
1756,47
1757,47
1758,47
1759,47
1760,47
1761,47
1762,47
1763,47
1764,47
1765,47
1766,47
1767,47
1768,47
1769,47
1770,47
1771,47
1772,47
1773,47
1774,47
1775,47
1776,48
1777,48
1778,48
1779,48
1780,48
1781,48
1782,48
1783,48
1784,48
1785,48
1786,48
1787,48
1788,48
1789,48
1790,48
1791,48
1792,48
1793,48
1794,48
1795,48
1796,48
1797,48
1798,48
1799,48
1800,48
1801,48
1802,48
1803,48
1804,48
1805,48
1806,48
1807,48
1808,48
1809,48
1810,48
1811,48
1812,48
1813,49
1814,49
1815,49
1816,49
1817,49
1818,49
1819,49
1820,49
1821,49
1822,49
1823,49
1824,49
1825,49
1826,49
1827,49
1828,49
1829,49
1830,49
1831,49
1832,49
1833,49
1834,49
1835,49
1836,49
1837,49
1838,49
1839,49
1840,49
1841,49
1842,49
1843,49
1844,49
1845,49
1846,49
1847,49
1848,49
1849,49
1850,50
1851,50
1852,50
1853,50
1854,50
1855,50
1856,50
1857,50
1858,50
1859,50
1860,50
1861,50
1862,50
1863,50
1864,50
1865,50
1866,50
1867,50
1868,50
1869,50
1870,50
1871,50
1872,50
1873,50
1874,50
1875,50
1876,50
1877,50
1878,50
1879,50
1880,50
1881,50
1882,50
1883,50
1884,50
1885,50
1886,50
1887,51
1888,51
1889,51
1890,51
1891,51
1892,51
1893,51
1894,51
1895,51
1896,51
1897,51
1898,51
1899,51
1900,51
1901,51
1902,51
1903,51
1904,51
1905,51
1906,51
1907,51
1908,51
1909,51
1910,51
1911,51
1912,51
1913,51
1914,51
1915,51
1916,51
1917,51
1918,51
1919,51
1920,51
1921,51
1922,51
1923,51
1924,52
1925,52
1926,52
1927,52
1928,52
1929,52
1930,52
1931,52
1932,52
1933,52
1934,52
1935,52
1936,52
1937,52
1938,52
1939,52
1940,52
1941,52
1942,52
1943,52
1944,52
1945,52
1946,52
1947,52
1948,52
1949,52
1950,52
1951,52
1952,52
1953,52
1954,52
1955,52
1956,52
1957,52
1958,52
1959,52
1960,52
1961,52
1962,53
1963,53
1964,53
1965,53
1966,53
1967,53
1968,53
1969,53
1970,53
1971,53
1972,53
1973,53
1974,53
1975,53
1976,53
1977,53
1978,53
1979,53
1980,53
1981,53
1982,53
1983,53
1984,53
1985,53
1986,53
1987,53
1988,53
1989,53
1990,53
1991,53
1992,53
1993,53
1994,53
1995,53
1996,53
1997,53
1998,53
1999,53
2000,54
2001,54
2002,54
2003,54
2004,54
2005,54
2006,54
2007,54
2008,54
2009,54
2010,54
2011,54
2012,54
2013,54
2014,54
2015,54
2016,54
2017,54
2018,54
2019,54
2020,54
2021,54
2022,54
2023,54
2024,54
2025,54
2026,54
2027,54
2028,54
2029,54
2030,54
2031,54
2032,54
2033,54
2034,54
2035,54
2036,54
2037,54
2038,55
2039,55
2040,55
2041,55
2042,55
2043,55
2044,55
2045,55
2046,55
2047,55
2048,55
2049,55
2050,55
2051,55
2052,55
2053,55
2054,55
2055,55
2056,55
2057,55
2058,55
2059,55
2060,55
2061,55
2062,55
2063,55
2064,55
2065,55
2066,55
2067,55
2068,55
2069,55
2070,55
2071,55
2072,55
2073,55
2074,55
2075,55
2076,56
2077,56
2078,56
2079,56
2080,56
2081,56
2082,56
2083,56
2084,56
2085,56
2086,56
2087,56
2088,56
2089,56
2090,56
2091,56
2092,56
2093,56
2094,56
2095,56
2096,56
2097,56
2098,56
2099,56
2100,56
2101,56
2102,56
2103,56
2104,56
2105,56
2106,56
2107,56
2108,56
2109,56
2110,56
2111,56
2112,56
2113,56
2114,57
2115,57
2116,57
2117,57
2118,57
2119,57
2120,57
2121,57
2122,57
2123,57
2124,57
2125,57
2126,57
2127,57
2128,57
2129,57
2130,57
2131,57
2132,57
2133,57
2134,57
2135,57
2136,57
2137,57
2138,57
2139,57
2140,57
2141,57
2142,57
2143,57
2144,57
2145,57
2146,57
2147,57
2148,57
2149,57
2150,57
2151,57
2152,58
2153,58
2154,58
2155,58
2156,58
2157,58
2158,58
2159,58
2160,58
2161,58
2162,58
2163,58
2164,58
2165,58
2166,58
2167,58
2168,58
2169,58
2170,58
2171,58
2172,58
2173,58
2174,58
2175,58
2176,58
2177,58
2178,58
2179,58
2180,58
2181,58
2182,58
2183,58
2184,58
2185,58
2186,58
2187,58
2188,58
2189,58
2190,59
2191,59
2192,59
2193,59
2194,59
2195,59
2196,59
2197,59
2198,59
2199,59
2200,59
2201,59
2202,59
2203,59
2204,59
2205,59
2206,59
2207,59
2208,59
2209,59
2210,59
2211,59
2212,59
2213,59
2214,59
2215,59
2216,59
2217,59
2218,59
2219,59
2220,59
2221,59
2222,59
2223,59
2224,59
2225,59
2226,59
2227,59
2228,60
2229,60
2230,60
2231,60
2232,60
2233,60
2234,60
2235,60
2236,60
2237,60
2238,60
2239,60
2240,60
2241,60
2242,60
2243,60
2244,60
2245,60
2246,60
2247,60
2248,60
2249,60
2250,60
2251,60
2252,60
2253,60
2254,60
2255,60
2256,60
2257,60
2258,60
2259,60
2260,60
2261,60
2262,60
2263,60
2264,60
2265,60
2266,61
2267,61
2268,61
2269,61
2270,61
2271,61
2272,61
2273,61
2274,61
2275,61
2276,61
2277,61
2278,61
2279,61
2280,61
2281,61
2282,61
2283,61
2284,61
2285,61
2286,61
2287,61
2288,61
2289,61
2290,61
2291,61
2292,61
2293,61
2294,61
2295,61
2296,61
2297,61
2298,61
2299,61
2300,61
2301,61
2302,61
2303,61
2304,62
2305,62
2306,62
2307,62
2308,62
2309,62
2310,62
2311,62
2312,62
2313,62
2314,62
2315,62
2316,62
2317,62
2318,62
2319,62
2320,62
2321,62
2322,62
2323,62
2324,62
2325,62
2326,62
2327,62
2328,62
2329,62
2330,62
2331,62
2332,62
2333,62
2334,62
2335,62
2336,62
2337,62
2338,62
2339,62
2340,62
2341,62
2342,63
2343,63
2344,63
2345,63
2346,63
2347,63
2348,63
2349,63
2350,63
2351,63
2352,63
2353,63
2354,63
2355,63
2356,63
2357,63
2358,63
2359,63
2360,63
2361,63
2362,63
2363,63
2364,63
2365,63
2366,63
2367,63
2368,63
2369,63
2370,63
2371,63
2372,63
2373,63
2374,63
2375,63
2376,63
2377,63
2378,63
2379,63
2380,64
2381,64
2382,64
2383,64
2384,64
2385,64
2386,64
2387,64
2388,64
2389,64
2390,64
2391,64
2392,64
2393,64
2394,64
2395,64
2396,64
2397,64
2398,64
2399,64
2400,64
2401,64
2402,64
2403,64
2404,64
2405,64
2406,64
2407,64
2408,64
2409,64
2410,64
2411,64
2412,64
2413,64
2414,64
2415,64
2416,64
2417,64
2418,65
2419,65
2420,65
2421,65
2422,65
2423,65
2424,65
2425,65
2426,65
2427,65
2428,65
2429,65
2430,65
2431,65
2432,65
2433,65
2434,65
2435,65
2436,65
2437,65
2438,65
2439,65
2440,65
2441,65
2442,65
2443,65
2444,65
2445,65
2446,65
2447,65
2448,65
2449,65
2450,65
2451,65
2452,65
2453,65
2454,65
2455,65
2456,66
2457,66
2458,66
2459,66
2460,66
2461,66
2462,66
2463,66
2464,66
2465,66
2466,66
2467,66
2468,66
2469,66
2470,66
2471,66
2472,66
2473,66
2474,66
2475,66
2476,66
2477,66
2478,66
2479,66
2480,66
2481,66
2482,66
2483,66
2484,66
2485,66
2486,66
2487,66
2488,66
2489,66
2490,66
2491,66
2492,66
2493,66
2494,67
2495,67
2496,67
2497,67
2498,67
2499,67
2500,67
2501,67
2502,67
2503,67
2504,67
2505,67
2506,67
2507,67
2508,67
2509,67
2510,67
2511,67
2512,67
2513,67
2514,67
2515,67
2516,67
2517,67
2518,67
2519,67
2520,67
2521,67
2522,67
2523,67
2524,67
2525,67
2526,67
2527,67
2528,67
2529,67
2530,67
2531,67
2532,68
2533,68
2534,68
2535,68
2536,68
2537,68
2538,68
2539,68
2540,68
2541,68
2542,68
2543,68
2544,68
2545,68
2546,68
2547,68
2548,68
2549,68
2550,68
2551,68
2552,68
2553,68
2554,68
2555,68
2556,68
2557,68
2558,68
2559,68
2560,68
2561,68
2562,68
2563,68
2564,68
2565,68
2566,68
2567,68
2568,68
2569,68
2570,69
2571,69
2572,69
2573,69
2574,69
2575,69
2576,69
2577,69
2578,69
2579,69
2580,69
2581,69
2582,69
2583,69
2584,69
2585,69
2586,69
2587,69
2588,69
2589,69
2590,69
2591,69
2592,69
2593,69
2594,69
2595,69
2596,69
2597,69
2598,69
2599,69
2600,69
2601,69
2602,69
2603,69
2604,69
2605,69
2606,69
2607,69
2608,70
2609,70
2610,70
2611,70
2612,70
2613,70
2614,70
2615,70
2616,70
2617,70
2618,70
2619,70
2620,70
2621,70
2622,70
2623,70
2624,70
2625,70
2626,70
2627,70
2628,70
2629,70
2630,70
2631,70
2632,70
2633,70
2634,70
2635,70
2636,70
2637,70
2638,70
2639,70
2640,70
2641,70
2642,70
2643,70
2644,70
2645,70
2646,71
2647,71
2648,71
2649,71
2650,71
2651,71
2652,71
2653,71
2654,71
2655,71
2656,71
2657,71
2658,71
2659,71
2660,71
2661,71
2662,71
2663,71
2664,71
2665,71
2666,71
2667,71
2668,71
2669,71
2670,71
2671,71
2672,71
2673,71
2674,71
2675,71
2676,71
2677,71
2678,71
2679,71
2680,71
2681,71
2682,71
2683,71
2684,72
2685,72
2686,72
2687,72
2688,72
2689,72
2690,72
2691,72
2692,72
2693,72
2694,72
2695,72
2696,72
2697,72
2698,72
2699,72
2700,72
2701,72
2702,72
2703,72
2704,72
2705,72
2706,72
2707,72
2708,72
2709,72
2710,72
2711,72
2712,72
2713,72
2714,72
2715,72
2716,72
2717,72
2718,72
2719,72
2720,72
2721,72
2722,73
2723,73
2724,73
2725,73
2726,73
2727,73
2728,73
2729,73
2730,73
2731,73
2732,73
2733,73
2734,73
2735,73
2736,73
2737,73
2738,73
2739,73
2740,73
2741,73
2742,73
2743,73
2744,73
2745,73
2746,73
2747,73
2748,73
2749,73
2750,73
2751,73
2752,73
2753,73
2754,73
2755,73
2756,73
2757,73
2758,73
2759,73
2760,74
2761,74
2762,74
2763,74
2764,74
2765,74
2766,74
2767,74
2768,74
2769,74
2770,74
2771,74
2772,74
2773,74
2774,74
2775,74
2776,74
2777,74
2778,74
2779,74
2780,74
2781,74
2782,74
2783,74
2784,74
2785,74
2786,74
2787,74
2788,74
2789,74
2790,74
2791,74
2792,74
2793,74
2794,74
2795,74
2796,74
2797,74
2798,75
2799,75
2800,75
2801,75
2802,75
2803,75
2804,75
2805,75
2806,75
2807,75
2808,75
2809,75
2810,75
2811,75
2812,75
2813,75
2814,75
2815,75
2816,75
2817,75
2818,75
2819,75
2820,75
2821,75
2822,75
2823,75
2824,75
2825,75
2826,75
2827,75
2828,75
2829,75
2830,75
2831,75
2832,75
2833,75
2834,75
2835,75
2836,76
2837,76
2838,76
2839,76
2840,76
2841,76
2842,76
2843,76
2844,76
2845,76
2846,76
2847,76
2848,76
2849,76
2850,76
2851,76
2852,76
2853,76
2854,76
2855,76
2856,76
2857,76
2858,76
2859,76
2860,76
2861,76
2862,76
2863,76
2864,76
2865,76
2866,76
2867,76
2868,76
2869,76
2870,76
2871,76
2872,76
2873,76
2874,77
2875,77
2876,77
2877,77
2878,77
2879,77
2880,77
2881,77
2882,77
2883,77
2884,77
2885,77
2886,77
2887,77
2888,77
2889,77
2890,77
2891,77
2892,77
2893,77
2894,77
2895,77
2896,77
2897,77
2898,77
2899,77
2900,77
2901,77
2902,77
2903,77
2904,77
2905,77
2906,77
2907,77
2908,77
2909,77
2910,77
2911,77
2912,78
2913,78
2914,78
2915,78
2916,78
2917,78
2918,78
2919,78
2920,78
2921,78
2922,78
2923,78
2924,78
2925,78
2926,78
2927,78
2928,78
2929,78
2930,78
2931,78
2932,78
2933,78
2934,78
2935,78
2936,78
2937,78
2938,78
2939,78
2940,78
2941,78
2942,78
2943,78
2944,78
2945,78
2946,78
2947,78
2948,78
2949,78
2950,79
2951,79
2952,79
2953,79
2954,79
2955,79
2956,79
2957,79
2958,79
2959,79
2960,79
2961,79
2962,79
2963,79
2964,79
2965,79
2966,79
2967,79
2968,79
2969,79
2970,79
2971,79
2972,79
2973,79
2974,79
2975,79
2976,79
2977,79
2978,79
2979,79
2980,79
2981,79
2982,79
2983,79
2984,79
2985,79
2986,79
2987,79
